�csaver
Saver
q )�q}q(X   dataq]q(}q(JR?�c__main__
User
q)�q}q(X   tg_idq	JR?�X   nameq
X   МаксимqX   roomqNX   wordsq]q(]q]q(X   аэропОртыqX
   бАнтыqX   бОродуqX   бухгАлтеровqX   вероисповЕданиеqX   граждАнствоqX
   дефИсqX   диспансЕрqX   договорЁнностьqX   докумЕнтqX
   досУгqX   еретИкqX   жалюзИqX   знАчимостьqX   ИксыqX   каталОгq X   монолОгq!X   квартАлq"X   киломЕтрq#X   кОнусыq$X   корЫстьq%X
   крАныq&X   кремЕньq'X   лЕкторыq(X
   лыжнЯq)X   мЕстностейq*X   мусоропровОдq+X   намЕрениеq,X   нарОстq-X   нЕдругq.X
   недУгq/X   некролОгq0X   нЕнавистьq1X   нОвостиq2X   нОготьq3X   Отрочествоq4X   партЕрq5X   портфЕльq6X   пОручниq7X   придАноеq8X   призЫвq9X
   отзЫвq:X   свЁклаq;X   сирОтыq<X   срЕдстваq=X
   созЫвq>X   столЯрq?X   тамОжняq@X
   тОртыqAX   цемЕнтqBX   цЕнтнерqCX   цепОчкаqDX
   шАрфыqEX
   шофЁрqFX   экспЕртqGX
   вернАqHX   красИвееqIX   красИвейшийqJX   кУхонныйqKX
   ловкАqLX   оптОвыйqMX   прозорлИваqNX   рядУqOX   болтлИваqPX   слИвовыйqQX   брАтьсяqRX   бралАсьqSX
   взятьqTX
   взялАqUX   взЯтьсяqVX   взялАсьqWX   включИтьqXX   включИшьqYX   включИтqZX   включИмq[X   влИтьсяq\X   влилАсьq]X   ворвАтьсяq^X   ворвалАсьq_X   воспринЯтьq`X   воспринялАqaX   воссоздАтьqbX   воссоздалАqcX   вручИтьqdX   вручИтqeX
   гнАтьqfX
   гналАqgX   гнАтьсяqhX   гналАсьqiX   добрАтьqjX   добралАqkX   добрАтьсяqlX   добралАсьqmX   дождАтьсяqnX   дождалАсьqoX   дозвонИтьсяqpX   дозвонИтсяqqX   дозвонЯтсяqrX   дозИроватьqsX
   ждатьqtX
   ждалАquX   жИтьсяqvX   жилОсьqwX   закУпоритьqxX   занЯтьqyX
   зАнялqzX   занялАq{X   зАнялоq|X   зАнялиq}X   заперЕтьq~X   заперлАqX   заперЕтьсяq�X   заперлАсьq�X
   зватьq�X
   звалАq�X   звонИтьq�X   звонИшьq�X   звонИтq�X   звонИмq�X   исчЕрпатьq�X
   клАлаq�X   клЕитьq�X   крАстьсяq�X   крАласьq�X
   лгатьq�X
   лгалАq�X   литьq�X   лилАq�X   лИтьсяq�X   лилАсьq�X   наврАтьq�X   наделИтьq�X   наделИтq�X   надорвАтьсяq�X   надорвалАсьq�X   назвАтьсяq�X   назвалАсьq�X   накренИтьсяq�X   накренИтсяq�X   налИтьq�X   налилАq�X   нарвАтьq�X   нарвалАq�X   насорИтьq�X   насорИтq�X   начАтьq�X
   нАчалq�X   началАq�X   нАчалиq�X   обзвонИтьq�X   обзвонИтq�X   облегчИтьq�X   облегчИтq�X   облИтьсяq�X   облилАсьq�X   обнЯтьсяq�X   обнялАсьq�X   обогнАтьq�X   обогналАq�X   ободрАтьq�X   ободралАq�X   ободрИтьq�X   ободрИтьсяq�X   ободрИшьсяq�X   обострИтьq�X   одолжИтq�X   озлОбитьq�X   оклЕитьq�X   окружИтьq�X   окружИтq�X   опломбировАтьq�X   формировАтьq�X   нормировАтьq�X   сортировАтьq�X   премировАтьq�X   опОшлитьq�X   освЕдомитьсяq�X   освЕдомишьсяq�X   отбЫтьq�X   отбылАq�X   отдАтьq�X   отдалАq�X   откУпоритьq�X   откУпорилq�X   отозвалАq�X   отозвАтьсяq�X   отозвалАсьq�X   перезвонИтьq�X   перезвонИтq�X   перелИтьq�X   перелилАq�X   плодоносИтьq�X   повторИтьq�X   повторИтq�X   позвАтьq�X   позвалАq�X   позвонИтьq�X   позвонИшьq�X   позвонИтq�X   полИтьq�X   полилАq�X   положИтьq�X   положИлq�X   понЯтьq�X   послАтьq�X   послАлаq�X   прибЫтьq�X   прИбылq�X   прибылАq�X   прИбылоq�X   принЯтьq�X   прИнялq�X   прИнялиq�X   принялАq�X   принУдитьq�X
   рвАтьq�X
   рвалАq�X   сверлИтьq�X   сверлИшьq�X   сверлИтq�X
   снЯтьq�X
   снялАq�X   создАтьq�X   создалАq�X   сорвАтьq�X   сорвалАq�X   сорИтьq�X
   сорИтq�X   убрАтьq�X   убралАq�X   убыстрИтьq�X   углубИтьq�X   укрепИтьq�X   укрепИтq�X   чЕрпатьq�X   щемИтьq�X
   щемИтq�X   щЁлкатьq�X   балОванныйq�X   включЁнныйr   X   включЁнr  X   низведЁнныйr  X   довезЁнныйr  X   зАгнутыйr  X   зАнятыйr  X   занятАr  X   зАпертыйr  X   заселЁнныйr  X   избалОванныйr	  X   балОванныйr
  X   кормЯщийr  X   кровоточАщийr  X   молЯщийr  X   нажИвшийr  X   нАжитыйr  X   нажитАr  X   налИвшийr  X   налитАr  X   нанЯвшийся	r  X   начАвшийr  X   нАчатыйr  X   низведЁнныйr  X   низведЁнr  X   включЁнныйr  X   ободрЁнныйr  X   ободрЁнr  X   ободренАr  X   обострЁнныйr  X   отключЁнныйr  X   определЁнныйr  X   определЁнr  X   отключЁнныйr   X   повторЁнныйr!  X   поделЁнныйr"  X   понЯвшийr#  X   прИнятыйr$  X   приручЁнныйr%  X   прожИвшийr&  X   снЯтыйr'  X
   снятАr(  X   сОгнутыйr)  X   балУясьr*  X   закУпоривr+  X
   начАвr,  X   начАвшисьr-  X   поднЯвr.  X
   понЯвr/  X   прибЫвr0  X   вОвремяr1  X   добелАr2  X   дОверхуr3  X   донЕльзяr4  X   дОсухаr5  X   завИдноr6  X   зАгодяr7  X   зАсветлоr8  X   зАтемноr9  X   красИвееr:  X   навЕрхr;  X   надОлгоr<  X   ненадОлгоr=  e]r>  eX   statsr?  }r@  (X   заселенАrA  ]rB  (KK K eX   одолжИтьrC  ]rD  (KK K eX   отозвАтьrE  ]rF  (KK K eX   клАстьrG  ]rH  (KK K eh�]rI  (KK KeX
   отдАвrJ  ]rK  (KK K ehJ]rL  (KK KeX   стАтуяrM  ]rN  (KK K eX   навралАrO  ]rP  (KK K eX   понялАrQ  ]rR  (KK K ej   ]rS  (KK Keh`]rT  (KK K eh�]rU  (KK Kehh]rV  (KK K ej  ]rW  (KK K eX   дОнизуrX  ]rY  (KK K eX   запертАrZ  ]r[  (KK K euX	   last_wordr\  h�X	   favouriter]  ]r^  h�aX
   prohibitedr_  ]r`  (jA  jC  jE  jG  jJ  jM  jO  jQ  jX  jZ  eubJ�]h)�ra  }rb  (h	J�]h
X   edombekrc  hNh]rd  (]re  ]rf  (X   аэропОртыrg  X
   бАнтыrh  X   бОродуri  X   бухгАлтеровrj  X   вероисповЕданиеrk  X   граждАнствоrl  X
   дефИсrm  X   диспансЕрrn  X   договорЁнностьro  X   докумЕнтrp  X
   досУгrq  X   еретИкrr  X   жалюзИrs  X   знАчимостьrt  X   Иксыru  X   каталОгrv  X   монолОгrw  X   квартАлrx  X   киломЕтрry  X   кОнусыrz  X   корЫстьr{  X
   крАныr|  X   кремЕньr}  X   лЕкторыr~  X
   лыжнЯr  X   мЕстностейr�  X   мусоропровОдr�  X   намЕрениеr�  X   нарОстr�  X   нЕдругr�  X
   недУгr�  X   некролОгr�  X   нЕнавистьr�  X   нОвостиr�  X   нОготьr�  X   Отрочествоr�  X   партЕрr�  X   портфЕльr�  X   пОручниr�  X   придАноеr�  X   призЫвr�  X
   отзЫвr�  X   свЁклаr�  X   сирОтыr�  X   срЕдстваr�  X
   созЫвr�  X   стАтуяr�  X   столЯрr�  X   тамОжняr�  X
   тОртыr�  X   цемЕнтr�  X   цЕнтнерr�  X   цепОчкаr�  X
   шАрфыr�  X
   шофЁрr�  X   экспЕртr�  X
   вернАr�  X   красИвееr�  X   красИвейшийr�  X   кУхонныйr�  X
   ловкАr�  X   оптОвыйr�  X   прозорлИваr�  X   рядУr�  X   болтлИваr�  X   слИвовыйr�  X   брАтьсяr�  X   бралАсьr�  X
   взятьr�  X
   взялАr�  X   взЯтьсяr�  X   взялАсьr�  X   включИтьr�  X   включИшьr�  X   включИтr�  X   включИмr�  X   влИтьсяr�  X   влилАсьr�  X   ворвАтьсяr�  X   ворвалАсьr�  X   воспринЯтьr�  X   воспринялАr�  X   воссоздАтьr�  X   воссоздалАr�  X   вручИтьr�  X   вручИтr�  X
   гнАтьr�  X
   гналАr�  X   гнАтьсяr�  X   гналАсьr�  X   добрАтьr�  X   добралАr�  X   добрАтьсяr�  X   добралАсьr�  X   дождАтьсяr�  X   дождалАсьr�  X   дозвонИтьсяr�  X   дозвонИтсяr�  X   дозвонЯтсяr�  X   дозИроватьr�  X
   ждатьr�  X
   ждалАr�  X   жИтьсяr�  X   жилОсьr�  X   закУпоритьr�  X   занЯтьr�  X
   зАнялr�  X   занялАr�  X   зАнялоr�  X   зАнялиr�  X   заперЕтьr�  X   заперлАr�  X   заперЕтьсяr�  X   заперлАсьr�  X
   зватьr�  X
   звалАr�  X   звонИтьr�  X   звонИшьr�  X   звонИтr�  X   звонИмr�  X   исчЕрпатьr�  X   клАстьr�  X
   клАлаr�  X   клЕитьr�  X   крАстьсяr�  X   крАласьr�  X
   лгатьr�  X
   лгалАr�  X   литьr�  X   лилАr�  X   лИтьсяr�  X   лилАсьr�  X   наврАтьr�  X   навралАr�  X   наделИтьr�  X   наделИтr�  X   надорвАтьсяr�  X   надорвалАсьr�  X   назвАтьсяr�  X   назвалАсьr�  X   накренИтьсяr�  X   накренИтсяr�  X   налИтьr�  X   нарвАтьr�  X   нарвалАr�  X   насорИтьr�  X   насорИтr�  X   начАтьr�  X
   нАчалr�  X   началАr�  X   нАчалиr�  X   обзвонИтьr�  X   обзвонИтr�  X   облегчИтьr   X   облегчИтr  X   облИтьсяr  X   облилАсьr  X   обнЯтьсяr  X   обнялАсьr  X   обогнАтьr  X   обогналАr  X   ободрАтьr  X   ободралАr	  X   ободрИтьr
  X   ободрИтьсяr  X   ободрИшьсяr  X   обострИтьr  X   одолжИтьr  X   одолжИтr  X   озлОбитьr  X   оклЕитьr  X   окружИтьr  X   окружИтr  X   опломбировАтьr  X   формировАтьr  X   нормировАтьr  X   сортировАтьr  X   премировАтьr  X   опОшлитьr  X   освЕдомитьсяr  X   освЕдомишьсяr  X   отбЫтьr  X   отбылАr  X   отдАтьr  X   отдалАr  X   откУпоритьr   X   откУпорилr!  X   отозвАтьr"  X   отозвалАr#  X   отозвАтьсяr$  X   отозвалАсьr%  X   перезвонИтьr&  X   перезвонИтr'  X   перелИтьr(  X   перелилАr)  X   плодоносИтьr*  X   повторИтьr+  X   повторИтr,  X   позвАтьr-  X   позвалАr.  X   позвонИтьr/  X   позвонИшьr0  X   позвонИтr1  X   полИтьr2  X   полилАr3  X   положИтьr4  X   положИлr5  X   понЯтьr6  X   понялАr7  X   послАтьr8  X   послАлаr9  X   прибЫтьr:  X   прИбылr;  X   прибылАr<  X   прИбылоr=  X   принЯтьr>  X   прИнялr?  X   прИнялиr@  X   принялАrA  X   принУдитьrB  X
   рвАтьrC  X
   рвалАrD  X   сверлИтьrE  X   сверлИшьrF  X   сверлИтrG  X
   снЯтьrH  X
   снялАrI  X   создАтьrJ  X   создалАrK  X   сорвАтьrL  X   сорвалАrM  X   сорИтьrN  X
   сорИтrO  X   убрАтьrP  X   убралАrQ  X   убыстрИтьrR  X   углубИтьrS  X   укрепИтьrT  X   укрепИтrU  X   чЕрпатьrV  X   щемИтьrW  X
   щемИтrX  X   щЁлкатьrY  X   балОванныйrZ  X   включЁнныйr[  X   включЁнr\  X   низведЁнныйr]  X   довезЁнныйr^  X   зАгнутыйr_  X   зАнятыйr`  X   занятАra  X   зАпертыйrb  X   запертАrc  X   заселЁнныйrd  X   заселенАre  X   избалОванныйrf  X   балОванныйrg  X   кормЯщийrh  X   кровоточАщийri  X   молЯщийrj  X   нажИвшийrk  X   нАжитыйrl  X   нажитАrm  X   налИвшийrn  X   налитАro  X   нанЯвшийся	rp  X   начАвшийrq  X   нАчатыйrr  X   низведЁнныйrs  X   низведЁнrt  X   включЁнныйru  X   ободрЁнныйrv  X   ободрЁнrw  X   ободренАrx  X   обострЁнныйry  X   отключЁнныйrz  X   определЁнныйr{  X   определЁнr|  X   отключЁнныйr}  X   повторЁнныйr~  X   поделЁнныйr  X   понЯвшийr�  X   прИнятыйr�  X   приручЁнныйr�  X   прожИвшийr�  X   снЯтыйr�  X
   снятАr�  X   сОгнутыйr�  X   балУясьr�  X   закУпоривr�  X
   начАвr�  X   начАвшисьr�  X
   отдАвr�  X   поднЯвr�  X
   понЯвr�  X   прибЫвr�  X   вОвремяr�  X   добелАr�  X   дОверхуr�  X   донЕльзяr�  X   дОнизуr�  X   дОсухаr�  X   завИдноr�  X   зАгодяr�  X   зАсветлоr�  X   зАтемноr�  X   красИвееr�  X   навЕрхr�  X   надОлгоr�  X   ненадОлгоr�  e]r�  ej?  }r�  (j  ]r�  (KK Kej  ]r�  (KK K ej  ]r�  (KK Kej�  ]r�  (KK KeX   налилАr�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (K KK ej�  ]r�  (KK K euj\  j5  j]  ]r�  j�  aj_  ]r�  j�  aubJ�&-h)�r�  }r�  (h	J�&-h
X   Александрr�  hNh]r�  (]r�  ]r�  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  (j>  ]r�  (K KKej�  ]r�  (KK Keuj\  j�  j]  ]r�  j_  ]r�  ubJ#J7%h)�r�  }r�  (h	J#J7%h
X   Glebr�  hNh]r�  (]r�  ]r�  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  j�  ]r�  (K KK esj\  j�  j]  ]r�  j�  aj_  ]r�  j�  aubJ���h)�r�  }r�  (h	J���h
X
   Антонr�  hNh]r�  (]r�  ]r�  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  (j=  ]r�  (KK Kej  ]r�  (KK K ej�  ]r�  (KK Keju  ]r�  (KK Kejn  ]r�  (KK K eja  ]r�  (KK Kej(  ]r�  (KK K ej�  ]r�  (KK K eji  ]r�  (KK K ejp  ]r�  (KK Kej|  ]r�  (KK K ej	  ]r�  (KK Keuj\  j�  j]  ]r�  j_  ]r�  ubJN<�!h)�r�  }r�  (h	JN<�!h
X   Marinar�  hNh]r�  (]r�  ]r�  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  j\  j  j]  ]r�  j_  ]r�  ubJl��!h)�r�  }r�  (h	Jl��!h
X   Машаr�  hNh]r�  (]r�  ]r�  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  (j�  ]r�  (KK K ejK  ]r�  (KK K ejR  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej=  ]r�  (KK K ej  ]r�  (K KKeuj\  j�  j]  ]r�  jK  aj_  ]r�  ubJ�<�.h)�r�  }r�  (h	J�<�.h
X   Polinar�  hNh]r�  (]r�  ]r�  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  (j1  ]r�  (KK K ej  ]r�  (KK K ejN  ]r   (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej  ]r  (KK K ejv  ]r  (KK K ejC  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ejy  ]r	  (KK K ejf  ]r
  (KK K ej  ]r  (KK K ej�  ]r  (KK K ejl  ]r  (K KKej�  ]r  (KK K ej�  ]r  (KK K ejM  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ejE  ]r  (KK K ej�  ]r  (KK K ejt  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ejs  ]r  (KK K ej�  ]r  (KK K ej  ]r  (KK K ej3  ]r  (KK K ej  ]r  (KK K ej)  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r   (KK K ej�  ]r!  (KK K ej;  ]r"  (KK K ej  ]r#  (KK K ej
  ]r$  (KK K ej�  ]r%  (KK K ej�  ]r&  (KK K ejP  ]r'  (KK K ej\  ]r(  (KK K ej�  ]r)  (KK K ej(  ]r*  (KK K ejF  ]r+  (KK K ej�  ]r,  (KK K ej�  ]r-  (KK K ej  ]r.  (KK K ej�  ]r/  (KK K ej�  ]r0  (KK K ej�  ]r1  (KK K ej  ]r2  (KK K ej�  ]r3  (KK K ej9  ]r4  (K KK euj\  j�  j]  ]r5  j_  ]r6  ubJ��-h)�r7  }r8  (h	J��-h
X   Васичекr9  hNh]r:  (]r;  ]r<  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r=  ej?  }r>  j\  j�  j]  ]r?  j_  ]r@  ubJ�Xl9h)�rA  }rB  (h	J�Xl9h
X   ВладиславrC  hNh]rD  (]rE  ]rF  (X   аэропОртыrG  X
   бАнтыrH  X   бОродуrI  X   бухгАлтеровrJ  X   вероисповЕданиеrK  X   граждАнствоrL  X
   дефИсrM  X   диспансЕрrN  X   договорЁнностьrO  X   докумЕнтrP  X
   досУгrQ  X   еретИкrR  X   жалюзИrS  X   знАчимостьrT  X   ИксыrU  X   каталОгrV  X   монолОгrW  X   квартАлrX  X   киломЕтрrY  X   кОнусыrZ  X   корЫстьr[  X
   крАныr\  X   кремЕньr]  X   лЕкторыr^  X
   лыжнЯr_  X   мЕстностейr`  X   мусоропровОдra  X   намЕрениеrb  X   нарОстrc  X   нЕдругrd  X
   недУгre  X   некролОгrf  X   нЕнавистьrg  X   нОвостиrh  X   нОготьri  X   Отрочествоrj  X   партЕрrk  X   портфЕльrl  X   пОручниrm  X   придАноеrn  X   призЫвro  X
   отзЫвrp  X   свЁклаrq  X   сирОтыrr  X   срЕдстваrs  X
   созЫвrt  X   стАтуяru  X   столЯрrv  X   тамОжняrw  X
   тОртыrx  X   цемЕнтry  X   цЕнтнерrz  X   цепОчкаr{  X
   шАрфыr|  X
   шофЁрr}  X   экспЕртr~  X
   вернАr  X   красИвееr�  X   красИвейшийr�  X   кУхонныйr�  X
   ловкАr�  X   оптОвыйr�  X   прозорлИваr�  X   рядУr�  X   болтлИваr�  X   слИвовыйr�  X   брАтьсяr�  X   бралАсьr�  X
   взятьr�  X
   взялАr�  X   взЯтьсяr�  X   взялАсьr�  X   включИтьr�  X   включИшьr�  X   включИтr�  X   включИмr�  X   влИтьсяr�  X   влилАсьr�  X   ворвАтьсяr�  X   ворвалАсьr�  X   воспринЯтьr�  X   воспринялАr�  X   воссоздАтьr�  X   воссоздалАr�  X   вручИтьr�  X   вручИтr�  X
   гнАтьr�  X
   гналАr�  X   гнАтьсяr�  X   гналАсьr�  X   добрАтьr�  X   добралАr�  X   добрАтьсяr�  X   добралАсьr�  X   дождАтьсяr�  X   дождалАсьr�  X   дозвонИтьсяr�  X   дозвонИтсяr�  X   дозвонЯтсяr�  X   дозИроватьr�  X
   ждатьr�  X
   ждалАr�  X   жИтьсяr�  X   жилОсьr�  X   закУпоритьr�  X   занЯтьr�  X
   зАнялr�  X   занялАr�  X   зАнялоr�  X   зАнялиr�  X   заперЕтьr�  X   заперлАr�  X   заперЕтьсяr�  X   заперлАсьr�  X
   зватьr�  X
   звалАr�  X   звонИтьr�  X   звонИшьr�  X   звонИтr�  X   звонИмr�  X   исчЕрпатьr�  X   клАстьr�  X
   клАлаr�  X   клЕитьr�  X   крАстьсяr�  X   крАласьr�  X
   лгалАr�  X   литьr�  X   лилАr�  X   лИтьсяr�  X   лилАсьr�  X   наврАтьr�  X   навралАr�  X   наделИтьr�  X   наделИтr�  X   надорвАтьсяr�  X   надорвалАсьr�  X   назвАтьсяr�  X   назвалАсьr�  X   накренИтьсяr�  X   накренИтсяr�  X   налИтьr�  X   налилАr�  X   нарвАтьr�  X   нарвалАr�  X   насорИтьr�  X   насорИтr�  X   начАтьr�  X
   нАчалr�  X   началАr�  X   нАчалиr�  X   обзвонИтьr�  X   обзвонИтr�  X   облегчИтьr�  X   облегчИтr�  X   облИтьсяr�  X   облилАсьr�  X   обнЯтьсяr�  X   обнялАсьr�  X   обогнАтьr�  X   обогналАr�  X   ободрАтьr�  X   ободралАr�  X   ободрИтьr�  X   ободрИтьсяr�  X   ободрИшьсяr�  X   обострИтьr�  X   одолжИтьr�  X   одолжИтr�  X   озлОбитьr�  X   оклЕитьr�  X   окружИтьr�  X   окружИтr�  X   опломбировАтьr�  X   формировАтьr�  X   нормировАтьr�  X   сортировАтьr�  X   премировАтьr�  X   опОшлитьr�  X   освЕдомитьсяr�  X   освЕдомишьсяr�  X   отбЫтьr�  X   отбылАr�  X   отдАтьr�  X   отдалАr�  X   откУпоритьr   X   откУпорилr  X   отозвАтьr  X   отозвалАr  X   отозвАтьсяr  X   отозвалАсьr  X   перезвонИтьr  X   перезвонИтr  X   перелИтьr  X   перелилАr	  X   плодоносИтьr
  X   повторИтьr  X   повторИтr  X   позвАтьr  X   позвалАr  X   позвонИтьr  X   позвонИшьr  X   позвонИтr  X   полИтьr  X   полилАr  X   положИтьr  X   положИлr  X   понЯтьr  X   понялАr  X   послАтьr  X   послАлаr  X   прибЫтьr  X   прИбылr  X   прибылАr  X   прИбылоr  X   принЯтьr  X   прИнялr  X   прИнялиr   X   принялАr!  X   принУдитьr"  X
   рвАтьr#  X
   рвалАr$  X   сверлИтьr%  X   сверлИшьr&  X   сверлИтr'  X
   снЯтьr(  X
   снялАr)  X   создАтьr*  X   создалАr+  X   сорвАтьr,  X   сорвалАr-  X   сорИтьr.  X
   сорИтr/  X   убрАтьr0  X   убралАr1  X   убыстрИтьr2  X   углубИтьr3  X   укрепИтьr4  X   укрепИтr5  X   чЕрпатьr6  X   щемИтьr7  X
   щемИтr8  X   щЁлкатьr9  X   балОванныйr:  X   включЁнныйr;  X   включЁнr<  X   низведЁнныйr=  X   довезЁнныйr>  X   зАгнутыйr?  X   зАнятыйr@  X   занятАrA  X   зАпертыйrB  X   запертАrC  X   заселЁнныйrD  X   заселенАrE  X   избалОванныйrF  X   балОванныйrG  X   кормЯщийrH  X   кровоточАщийrI  X   молЯщийrJ  X   нажИвшийrK  X   нАжитыйrL  X   нажитАrM  X   налИвшийrN  X   налитАrO  X   нанЯвшийся	rP  X   начАвшийrQ  X   нАчатыйrR  X   низведЁнныйrS  X   низведЁнrT  X   включЁнныйrU  X   ободрЁнныйrV  X   ободрЁнrW  X   ободренАrX  X   обострЁнныйrY  X   отключЁнныйrZ  X   определЁнныйr[  X   определЁнr\  X   отключЁнныйr]  X   повторЁнныйr^  X   поделЁнныйr_  X   понЯвшийr`  X   прИнятыйra  X   приручЁнныйrb  X   прожИвшийrc  X   снЯтыйrd  X
   снятАre  X   сОгнутыйrf  X   балУясьrg  X   закУпоривrh  X
   начАвri  X   начАвшисьrj  X
   отдАвrk  X   поднЯвrl  X
   понЯвrm  X   прибЫвrn  X   вОвремяro  X   добелАrp  X   дОверхуrq  X   донЕльзяrr  X   дОнизуrs  X   дОсухаrt  X   завИдноru  X   зАгодяrv  X   зАсветлоrw  X   зАтемноrx  X   красИвееry  X   навЕрхrz  X   надОлгоr{  X   ненадОлгоr|  e]r}  ej?  }r~  (ji  ]r  (KK Kej�  ]r�  (KK Kej  ]r�  (KK Kej/  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK Kej8  ]r�  (KK KeX
   лгатьr�  ]r�  (KK Kejj  ]r�  (KK Kej�  ]r�  (KK K ejP  ]r�  (KK Kej?  ]r�  (KK K ej"  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KKKejC  ]r�  (KK Kej�  ]r�  (KK Kej'  ]r�  (KK Kej[  ]r�  (KK KejY  ]r�  (KK Kej�  ]r�  (K KKejO  ]r�  (K KKej>  ]r�  (K KKej  ]r�  (K KKeuj\  j�  j]  ]r�  (ji  j�  ej_  ]r�  j�  aubJlz0"h)�r�  }r�  (h	Jlz0"h
X   Ikitr�  hNh]r�  (]r�  ]r�  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  (jE  ]r�  (KK K ejk  ]r�  (KK K ejs  ]r�  (KK K ej�  ]r�  (KK K ejj  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (K KK ej%  ]r�  (KK K ej�  ]r�  (KK K ejf  ]r�  (KK K ejp  ]r�  (KK K ej  ]r�  (KK K ejL  ]r�  (KK K ejg  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejd  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (K KKej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej}  ]r�  (KK K ej\  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej_  ]r�  (KK K ej  ]r�  (KK K ejD  ]r�  (KK K ej.  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejS  ]r�  (KK K ej�  ]r�  (KK K ejm  ]r�  (KK K ej
  ]r�  (KK K ej  ]r�  (KK K ej  ]r�  (KK K ej@  ]r�  (KK K ej  ]r�  (KK K ejj  ]r�  (KK K ej�  ]r�  (KK K ej3  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej{  ]r�  (KK K ejM  ]r�  (KK K ej�  ]r�  (KK K ej*  ]r�  (KK K eji  ]r�  (KK K ej�  ]r�  (KK K ej+  ]r�  (KK K ej�  ]r�  (KK K ej;  ]r�  (KK KejR  ]r�  (KK K ej2  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K eju  ]r�  (KK K ej>  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejC  ]r�  (KK K ejY  ]r�  (K KKej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejU  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K euj\  j�  j]  ]r�  j_  ]r�  ubJ�?�h)�r�  }r�  (h	J�?�h
X
   Борисr   hNh]r  (]r  ]r  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r  ej?  }r  (j�  ]r  (KK KejB  ]r  (KK Kej1  ]r  (KK K ej�  ]r	  (KK K ej�  ]r
  (KK K ej�  ]r  (KK K ejr  ]r  (KK K ej4  ]r  (KK K ejS  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej  ]r  (KK K ej�  ]r  (KK K ejo  ]r  (KK K ej  ]r  (KK KejA  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej{  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ejc  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej  ]r   (KK K ejW  ]r!  (KK Keuj\  j�  j]  ]r"  j_  ]r#  (j�  jc  j�  j  eubJ��_#h)�r$  }r%  (h	J��_#h
X   Степанr&  hNh]r'  (]r(  ]r)  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r*  ej?  }r+  (j   ]r,  (KK Kej�  ]r-  (KK Kej�  ]r.  (KK Kejr  ]r/  (KK Kej�  ]r0  (KK Kejc  ]r1  (KK Kej�  ]r2  (KK Kejs  ]r3  (K KKej�  ]r4  (KK Kej0  ]r5  (KK Kej�  ]r6  (KK Kej[  ]r7  (KK Kej  ]r8  (KK Kej�  ]r9  (KK Kej1  ]r:  (KK Kej�  ]r;  (KK Kej\  ]r<  (KK Kej�  ]r=  (KK Kej�  ]r>  (K KKej  ]r?  (KK Keuj\  j�  j]  ]r@  j_  ]rA  ubJ��h)�rB  }rC  (h	J��h
X   Lil telegramrD  hNh]rE  (]rF  ]rG  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]rH  ej?  }rI  (j�  ]rJ  (KK K ej�  ]rK  (KK K ejs  ]rL  (KK K ej�  ]rM  (KK K ejd  ]rN  (KK K ej  ]rO  (KK K ej�  ]rP  (KK K ej<  ]rQ  (KK K ej�  ]rR  (KK K ej�  ]rS  (KK K ej�  ]rT  (KK K ej�  ]rU  (KK K ej�  ]rV  (KK K euj\  j�  j]  ]rW  j_  ]rX  ubJos�h)�rY  }rZ  (h	Jos�h
X   Alinar[  hNh]r\  (]r]  ]r^  (jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r_  ej?  }r`  (j~  ]ra  (KK K ejh  ]rb  (KK K ej�  ]rc  (KK K ejk  ]rd  (KK K ej�  ]re  (KK K ej{  ]rf  (KK K ej�  ]rg  (K KKej�  ]rh  (KK K ej|  ]ri  (KK K ej�  ]rj  (KK K ej�  ]rk  (KK K ej.  ]rl  (KK K ej�  ]rm  (K KKej  ]rn  (KK K ejc  ]ro  (KK K ej�  ]rp  (KK K ej�  ]rq  (KK K ej�  ]rr  (KK K ejr  ]rs  (K KKej�  ]rt  (KK K ejA  ]ru  (KK K ej�  ]rv  (KK K ej�  ]rw  (KK K ej�  ]rx  (KK K ejM  ]ry  (KK K ej�  ]rz  (KK K ej�  ]r{  (KK K ej6  ]r|  (KK K ej�  ]r}  (KK K ej�  ]r~  (KK K ej'  ]r  (KK K ej�  ]r�  (KK K ejl  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej3  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej,  ]r�  (KK K ej�  ]r�  (KK K ejy  ]r�  (KK K ej�  ]r�  (KK K euj\  j�  j]  ]r�  j_  ]r�  ubJ���5h)�r�  }r�  (h	J���5h
X   Сергейr�  hNh]r�  (]r�  ]r�  (X   аэропОртыr�  X
   бАнтыr�  X   бОродуr�  X   бухгАлтеровr�  X   вероисповЕданиеr�  X   граждАнствоr�  X
   дефИсr�  X   диспансЕрr�  X   договорЁнностьr�  X   докумЕнтr�  X
   досУгr�  X   еретИкr�  X   жалюзИr�  X   знАчимостьr�  X   Иксыr�  X   каталОгr�  X   монолОгr�  X   квартАлr�  X   киломЕтрr�  X   кОнусыr�  X   корЫстьr�  X
   крАныr�  X   кремЕньr�  X   лЕкторыr�  X
   лыжнЯr�  X   мЕстностейr�  X   мусоропровОдr�  X   намЕрениеr�  X   нарОстr�  X   нЕдругr�  X
   недУгr�  X   некролОгr�  X   нЕнавистьr�  X   нОвостиr�  X   нОготьr�  X   Отрочествоr�  X   партЕрr�  X   портфЕльr�  X   пОручниr�  X   придАноеr�  X   призЫвr�  X
   отзЫвr�  X   свЁклаr�  X   сирОтыr�  X   срЕдстваr�  X
   созЫвr�  X   стАтуяr�  X   столЯрr�  X   тамОжняr�  X
   тОртыr�  X   цемЕнтr�  X   цЕнтнерr�  X   цепОчкаr�  X
   шАрфыr�  X
   шофЁрr�  X   экспЕртr�  X
   вернАr�  X   красИвееr�  X   красИвейшийr�  X   кУхонныйr�  X
   ловкАr�  X   оптОвыйr�  X   прозорлИваr�  X   рядУr�  X   болтлИваr�  X   слИвовыйr�  X   брАтьсяr�  X   бралАсьr�  X
   взятьr�  X
   взялАr�  X   взЯтьсяr�  X   взялАсьr�  X   включИтьr�  X   включИшьr�  X   включИтr�  X   включИмr�  X   влИтьсяr�  X   влилАсьr�  X   ворвАтьсяr�  X   ворвалАсьr�  X   воспринЯтьr�  X   воспринялАr�  X   воссоздАтьr�  X   воссоздалАr�  X   вручИтьr�  X   вручИтr�  X
   гнАтьr�  X
   гналАr�  X   гнАтьсяr�  X   гналАсьr�  X   добрАтьr�  X   добралАr�  X   добрАтьсяr�  X   добралАсьr�  X   дождАтьсяr�  X   дождалАсьr�  X   дозвонИтьсяr�  X   дозвонИтсяr�  X   дозвонЯтсяr�  X   дозИроватьr�  X
   ждатьr�  X
   ждалАr�  X   жИтьсяr�  X   жилОсьr�  X   закУпоритьr�  X   занЯтьr�  X
   зАнялr�  X   занялАr�  X   зАнялоr   X   зАнялиr  X   заперЕтьr  X   заперлАr  X   заперЕтьсяr  X   заперлАсьr  X
   зватьr  X
   звалАr  X   звонИтьr  X   звонИшьr	  X   звонИтr
  X   звонИмr  X   исчЕрпатьr  X   клАстьr  X
   клАлаr  X   клЕитьr  X   крАстьсяr  X   крАласьr  X
   лгатьr  X
   лгалАr  X   литьr  X   лилАr  X   лИтьсяr  X   лилАсьr  X   наврАтьr  X   навралАr  X   наделИтьr  X   наделИтr  X   надорвАтьсяr  X   надорвалАсьr  X   назвАтьсяr  X   назвалАсьr  X   накренИтьсяr   X   накренИтсяr!  X   налИтьr"  X   налилАr#  X   нарвАтьr$  X   нарвалАr%  X   насорИтьr&  X   насорИтr'  X   начАтьr(  X
   нАчалr)  X   началАr*  X   нАчалиr+  X   обзвонИтьr,  X   обзвонИтr-  X   облегчИтьr.  X   облегчИтr/  X   облИтьсяr0  X   облилАсьr1  X   обнЯтьсяr2  X   обнялАсьr3  X   обогнАтьr4  X   обогналАr5  X   ободрАтьr6  X   ободралАr7  X   ободрИтьr8  X   ободрИтьсяr9  X   ободрИшьсяr:  X   обострИтьr;  X   одолжИтьr<  X   одолжИтr=  X   озлОбитьr>  X   оклЕитьr?  X   окружИтьr@  X   окружИтrA  X   опломбировАтьrB  X   формировАтьrC  X   нормировАтьrD  X   сортировАтьrE  X   премировАтьrF  X   опОшлитьrG  X   освЕдомитьсяrH  X   освЕдомишьсяrI  X   отбЫтьrJ  X   отбылАrK  X   отдАтьrL  X   отдалАrM  X   откУпоритьrN  X   откУпорилrO  X   отозвАтьrP  X   отозвалАrQ  X   отозвАтьсяrR  X   отозвалАсьrS  X   перезвонИтьrT  X   перезвонИтrU  X   перелИтьrV  X   перелилАrW  X   плодоносИтьrX  X   повторИтьrY  X   повторИтrZ  X   позвАтьr[  X   позвалАr\  X   позвонИтьr]  X   позвонИшьr^  X   позвонИтr_  X   полИтьr`  X   полилАra  X   положИтьrb  X   положИлrc  X   понЯтьrd  X   понялАre  X   послАтьrf  X   послАлаrg  X   прибЫтьrh  X   прИбылri  X   прибылАrj  X   прИбылоrk  X   принЯтьrl  X   прИнялrm  X   прИнялиrn  X   принялАro  X   принУдитьrp  X
   рвАтьrq  X
   рвалАrr  X   сверлИтьrs  X   сверлИшьrt  X   сверлИтru  X
   снЯтьrv  X
   снялАrw  X   создАтьrx  X   создалАry  X   сорвАтьrz  X   сорвалАr{  X   сорИтьr|  X
   сорИтr}  X   убрАтьr~  X   убралАr  X   убыстрИтьr�  X   углубИтьr�  X   укрепИтьr�  X   укрепИтr�  X   чЕрпатьr�  X   щемИтьr�  X
   щемИтr�  X   щЁлкатьr�  X   балОванныйr�  X   включЁнныйr�  X   включЁнr�  X   низведЁнныйr�  X   довезЁнныйr�  X   зАгнутыйr�  X   зАнятыйr�  X   занятАr�  X   зАпертыйr�  X   запертАr�  X   заселЁнныйr�  X   заселенАr�  X   избалОванныйr�  X   балОванныйr�  X   кормЯщийr�  X   кровоточАщийr�  X   молЯщийr�  X   нажИвшийr�  X   нАжитыйr�  X   нажитАr�  X   налИвшийr�  X   налитАr�  X   нанЯвшийся	r�  X   начАвшийr�  X   нАчатыйr�  X   низведЁнныйr�  X   низведЁнr�  X   включЁнныйr�  X   ободрЁнныйr�  X   ободрЁнr�  X   ободренАr�  X   обострЁнныйr�  X   отключЁнныйr�  X   определЁнныйr�  X   определЁнr�  X   отключЁнныйr�  X   повторЁнныйr�  X   поделЁнныйr�  X   понЯвшийr�  X   прИнятыйr�  X   приручЁнныйr�  X   прожИвшийr�  X   снЯтыйr�  X
   снятАr�  X   сОгнутыйr�  X   балУясьr�  X   закУпоривr�  X
   начАвr�  X   начАвшисьr�  X
   отдАвr�  X   поднЯвr�  X
   понЯвr�  X   прибЫвr�  X   вОвремяr�  X   добелАr�  X   дОверхуr�  X   донЕльзяr�  X   дОнизуr�  X   дОсухаr�  X   завИдноr�  X   зАгодяr�  X   зАсветлоr�  X   зАтемноr�  X   красИвееr�  X   навЕрхr�  X   надОлгоr�  X   ненадОлгоr�  e]r�  ej?  }r�  (j�  ]r�  (KK K ej'  ]r�  (K KKej�  ]r�  (KK Kej\  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ejc  ]r�  (KK Kej�  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK K ej9  ]r�  (KK Keuj\  j�  j]  ]r�  j_  ]r�  ubJ5w�h)�r�  }r�  (h	J5w�h
X   Mumble Wizardr�  hNh]r�  (]r�  ]r�  (X   аэропОртыr�  X
   бАнтыr�  X   бОродуr�  X   бухгАлтеровr�  X   вероисповЕданиеr�  X   граждАнствоr�  X
   дефИсr�  X   диспансЕрr�  X   договорЁнностьr�  X   докумЕнтr�  X
   досУгr�  X   еретИкr�  X   жалюзИr�  X   знАчимостьr�  X   Иксыr�  X   каталОгr�  X   монолОгr�  X   квартАлr�  X   киломЕтрr�  X   кОнусыr�  X   корЫстьr�  X
   крАныr�  X   кремЕньr�  X   лЕкторыr�  X
   лыжнЯr�  X   мЕстностейr�  X   мусоропровОдr�  X   намЕрениеr�  X   нарОстr�  X   нЕдругr�  X
   недУгr   X   некролОгr  X   нЕнавистьr  X   нОвостиr  X   нОготьr  X   Отрочествоr  X   партЕрr  X   портфЕльr  X   пОручниr  X   придАноеr	  X   призЫвr
  X
   отзЫвr  X   свЁклаr  X   сирОтыr  X   срЕдстваr  X
   созЫвr  X   стАтуяr  X   столЯрr  X   тамОжняr  X
   тОртыr  X   цемЕнтr  X   цЕнтнерr  X   цепОчкаr  X
   шАрфыr  X
   шофЁрr  X   экспЕртr  X
   вернАr  X   красИвееr  X   красИвейшийr  X   кУхонныйr  X
   ловкАr  X   оптОвыйr  X   прозорлИваr   X   рядУr!  X   болтлИваr"  X   слИвовыйr#  X   брАтьсяr$  X   бралАсьr%  X
   взятьr&  X
   взялАr'  X   взЯтьсяr(  X   взялАсьr)  X   включИтьr*  X   включИшьr+  X   включИтr,  X   включИмr-  X   влИтьсяr.  X   влилАсьr/  X   ворвАтьсяr0  X   ворвалАсьr1  X   воспринЯтьr2  X   воспринялАr3  X   воссоздАтьr4  X   воссоздалАr5  X   вручИтьr6  X   вручИтr7  X
   гнАтьr8  X
   гналАr9  X   гнАтьсяr:  X   гналАсьr;  X   добрАтьr<  X   добралАr=  X   добрАтьсяr>  X   добралАсьr?  X   дождАтьсяr@  X   дождалАсьrA  X   дозвонИтьсяrB  X   дозвонИтсяrC  X   дозвонЯтсяrD  X   дозИроватьrE  X
   ждатьrF  X
   ждалАrG  X   жИтьсяrH  X   жилОсьrI  X   закУпоритьrJ  X   занЯтьrK  X
   зАнялrL  X   занялАrM  X   зАнялоrN  X   зАнялиrO  X   заперЕтьrP  X   заперлАrQ  X   заперЕтьсяrR  X   заперлАсьrS  X
   зватьrT  X
   звалАrU  X   звонИтьrV  X   звонИшьrW  X   звонИтrX  X   звонИмrY  X   исчЕрпатьrZ  X   клАстьr[  X
   клАлаr\  X   клЕитьr]  X   крАстьсяr^  X   крАласьr_  X
   лгатьr`  X
   лгалАra  X   литьrb  X   лилАrc  X   лИтьсяrd  X   лилАсьre  X   наврАтьrf  X   навралАrg  X   наделИтьrh  X   наделИтri  X   надорвАтьсяrj  X   надорвалАсьrk  X   назвАтьсяrl  X   назвалАсьrm  X   накренИтьсяrn  X   накренИтсяro  X   налИтьrp  X   налилАrq  X   нарвАтьrr  X   нарвалАrs  X   насорИтьrt  X   насорИтru  X   начАтьrv  X
   нАчалrw  X   началАrx  X   нАчалиry  X   обзвонИтьrz  X   обзвонИтr{  X   облегчИтьr|  X   облегчИтr}  X   облИтьсяr~  X   облилАсьr  X   обнЯтьсяr�  X   обнялАсьr�  X   обогнАтьr�  X   обогналАr�  X   ободрАтьr�  X   ободралАr�  X   ободрИтьr�  X   ободрИтьсяr�  X   ободрИшьсяr�  X   обострИтьr�  X   одолжИтьr�  X   одолжИтr�  X   озлОбитьr�  X   оклЕитьr�  X   окружИтьr�  X   окружИтr�  X   опломбировАтьr�  X   формировАтьr�  X   нормировАтьr�  X   сортировАтьr�  X   премировАтьr�  X   опОшлитьr�  X   освЕдомитьсяr�  X   освЕдомишьсяr�  X   отбЫтьr�  X   отбылАr�  X   отдАтьr�  X   отдалАr�  X   откУпоритьr�  X   откУпорилr�  X   отозвАтьr�  X   отозвалАr�  X   отозвАтьсяr�  X   отозвалАсьr�  X   перезвонИтьr�  X   перезвонИтr�  X   перелИтьr�  X   перелилАr�  X   плодоносИтьr�  X   повторИтьr�  X   повторИтr�  X   позвАтьr�  X   позвалАr�  X   позвонИтьr�  X   позвонИшьr�  X   позвонИтr�  X   полИтьr�  X   полилАr�  X   положИтьr�  X   положИлr�  X   понЯтьr�  X   понялАr�  X   послАтьr�  X   послАлаr�  X   прибЫтьr�  X   прИбылr�  X   прибылАr�  X   прИбылоr�  X   принЯтьr�  X   прИнялr�  X   прИнялиr�  X   принялАr�  X   принУдитьr�  X
   рвАтьr�  X
   рвалАr�  X   сверлИтьr�  X   сверлИшьr�  X   сверлИтr�  X
   снЯтьr�  X
   снялАr�  X   создАтьr�  X   создалАr�  X   сорвАтьr�  X   сорвалАr�  X   сорИтьr�  X
   сорИтr�  X   убрАтьr�  X   убралАr�  X   убыстрИтьr�  X   углубИтьr�  X   укрепИтьr�  X   укрепИтr�  X   чЕрпатьr�  X   щемИтьr�  X
   щемИтr�  X   щЁлкатьr�  X   балОванныйr�  X   включЁнныйr�  X   включЁнr�  X   низведЁнныйr�  X   довезЁнныйr�  X   зАгнутыйr�  X   зАнятыйr�  X   занятАr�  X   зАпертыйr�  X   запертАr�  X   заселЁнныйr�  X   заселенАr�  X   избалОванныйr�  X   балОванныйr�  X   кормЯщийr�  X   кровоточАщийr�  X   молЯщийr�  X   нажИвшийr�  X   нАжитыйr�  X   нажитАr�  X   налИвшийr�  X   налитАr�  X   нанЯвшийся	r�  X   начАвшийr�  X   нАчатыйr�  X   низведЁнныйr�  X   низведЁнr�  X   включЁнныйr�  X   ободрЁнныйr�  X   ободрЁнr�  X   ободренАr�  X   обострЁнныйr�  X   отключЁнныйr�  X   определЁнныйr�  X   определЁнr�  X   отключЁнныйr�  X   повторЁнныйr�  X   поделЁнныйr�  X   понЯвшийr�  X   прИнятыйr�  X   приручЁнныйr�  X   прожИвшийr�  X   снЯтыйr   X
   снятАr  X   сОгнутыйr  X   балУясьr  X   закУпоривr  X
   начАвr  X   начАвшисьr  X
   отдАвr  X   поднЯвr  X
   понЯвr	  X   прибЫвr
  X   вОвремяr  X   добелАr  X   дОверхуr  X   донЕльзяr  X   дОнизуr  X   дОсухаr  X   завИдноr  X   зАгодяr  X   зАсветлоr  X   зАтемноr  X   красИвееr  X   навЕрхr  X   надОлгоr  X   ненадОлгоr  e]r  ej?  }r  j\  j  j]  ]r  j_  ]r  ubJT�(h)�r  }r  (h	JT�(h
X   Mariar  hNh]r   (]r!  ]r"  (j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  e]r#  ej?  }r$  j\  j�  j]  ]r%  j_  ]r&  ubJbS�h)�r'  }r(  (h	JbS�h
X
   Иринаr)  hNh]r*  (]r+  ]r,  (hhhhhhhhhhhhhhhh h!h"h#h$h%h&h'h(h)h*h+h,h-h.h/h0h1h2h3h4h5h6h7h8h9h:h;h<h=h>jM  h?h@hAhBhChDhEhFhGhHhIhJhKhLhMhNhOhPhQhRhShThUhVhWhXhYhZh[h\h]h^h_h`hahbhchdhehfhghhhihjhkhlhmhnhohphqhrhshthuhvhwhxhyhzh{h|h}h~hh�h�h�h�h�h�h�h�h�jG  h�h�h�h�h�h�h�h�h�h�h�jO  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jC  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jE  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jQ  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�j   j  j  j  j  j  j  j  jZ  j  jA  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  jJ  j.  j/  j0  j1  j2  j3  j4  jX  j5  j6  j7  j8  j9  j:  j;  j<  j=  e]r-  ej?  }r.  (j  ]r/  (KK K ehr]r0  (KK K ej#  ]r1  (KK K ej.  ]r2  (KK K ehQ]r3  (KK Kej  ]r4  (KK Keh�]r5  (KK K ej  ]r6  (KK KehY]r7  (KK Kej;  ]r8  (KK K ejZ  ]r9  (KK K ehp]r:  (KK K ehM]r;  (KK K ehA]r<  (KK K eh*]r=  (KK K eh�]r>  (KK K eh^]r?  (KK K eh�]r@  (KK K eh�]rA  (KK K eh�]rB  (KK Keh�]rC  (KK K eh�]rD  (KK K eh�]rE  (KK K ehq]rF  (KK K eh�]rG  (KK K ehe]rH  (KK K eh>]rI  (KK K eh�]rJ  (KK K ej  ]rK  (KK K eh�]rL  (KK Kej  ]rM  (KK K eh�]rN  (KK K ej  ]rO  (KK K ej  ]rP  (KK K eh�]rQ  (KK Keh�]rR  (KK K eh�]rS  (KK K ehw]rT  (KK K eh�]rU  (KK K ejJ  ]rV  (KK K eh1]rW  (KK K ej<  ]rX  (KK K ejO  ]rY  (KK K eh�]rZ  (KK K eh�]r[  (KK K eh�]r\  (KK KejX  ]r]  (KK K ej+  ]r^  (KK K eh�]r_  (KK K ehI]r`  (KK K eh�]ra  (KK K eh�]rb  (KK K eh&]rc  (KK K eh�]rd  (KK K ej$  ]re  (KK K eh�]rf  (KK K ej   ]rg  (KK K eh]rh  (KK K eh8]ri  (KK K eh�]rj  (KK K ej  ]rk  (KK K eh]rl  (KK K eh6]rm  (KK K eh\]rn  (KK K eh%]ro  (KK K ehm]rp  (KK K eh�]rq  (KK K eh�]rr  (KK Keh]rs  (KK K ehf]rt  (KK K eh�]ru  (KK Keh]rv  (KK K ej  ]rw  (KK K ehP]rx  (KK K ej(  ]ry  (KK K eh�]rz  (KK K eh�]r{  (KK K eh�]r|  (KK K eh�]r}  (KK K eh_]r~  (KK K eh]r  (KK K eh�]r�  (KK K ej1  ]r�  (KK K eh�]r�  (KK K eh]r�  (KK K eh�]r�  (KK K eh�]r�  (KK K ehd]r�  (KK Keh�]r�  (KK K ehg]r�  (KK K eh�]r�  (KK K ejQ  ]r�  (KK K eh�]r�  (KK Keh�]r�  (KK K eh�]r�  (KK K eh�]r�  (KK K eh�]r�  (KKKeh�]r�  (KK K ej/  ]r�  (KK K ej	  ]r�  (KK K eh�]r�  (KK K eh]r�  (KK K ej  ]r�  (KK Keh�]r�  (KK K eh�]r�  (KK K euj\  jG  j]  ]r�  j_  ]r�  ubJ��f7h)�r�  }r�  (h	J��f7h
X   Катяr�  hNh]r�  (]r�  ]r�  (hhhhhhhhhhhhhhhh h!h"h#h$h%h&h'h(h)h*h+h,h-h.h/h0h1h2h3h4h5h6h7h8h9h:h;h<h=h>jM  h?h@hAhBhChDhEhFhGhHhIhJhKhLhMhNhOhPhQhRhShThUhVhWhXhYhZh[h\h]h^h_h`hahbhchdhehfhghhhihjhkhlhmhnhohphqhrhshthuhvhwhxhyhzh{h|h}h~hh�h�h�h�h�h�h�h�h�jG  h�h�h�h�h�h�h�h�h�h�h�jO  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jC  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jE  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jQ  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�j   j  j  j  j  j  j  j  jZ  j  jA  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  jJ  j.  j/  j0  j1  j2  j3  j4  jX  j5  j6  j7  j8  j9  j:  j;  j<  j=  e]r�  ej?  }r�  j\  h�j]  ]r�  j_  ]r�  ubJ1AN(h)�r�  }r�  (h	J1AN(h
X   Sashashr�  hNh]r�  (]r�  ]r�  (hhhhhhhhhhhhhhhh h!h"h#h$h%h&h'h(h)h*h+h,h-h.h/h0h1h2h3h4h5h6h7h8h9h:h;h<h=h>jM  h?h@hAhBhChDhEhFhGhHhIhJhKhLhMhNhOhPhQhRhShThUhVhWhXhYhZh[h\h]h^h_h`hahbhchdhehfhghhhihjhkhlhmhnhohphqhrhshthuhvhwhxhyhzh{h|h}h~hh�h�h�h�h�h�h�h�h�jG  h�h�h�h�h�h�h�h�h�h�h�jO  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jC  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jE  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�jQ  h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�h�j   j  j  j  j  j  j  j  jZ  j  jA  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  jJ  j.  j/  j0  j1  j2  j3  j4  jX  j5  j6  j7  j8  j9  j:  j;  j<  j=  e]r�  ej?  }r�  (hh]r�  (KK K ehL]r�  (KK K eh�]r�  (KK Kej(  ]r�  (KK K ej:  ]r�  (KK Keh�]r�  (K KKej  ]r�  (KK Keh]r�  (K KKeh,]r�  (KK K eh�]r�  (K KKeh�]r�  (K KKeh�]r�  (KK K eh�]r�  (KK K ehy]r�  (KK K eh�]r�  (KK K ej  ]r�  (KK K ehT]r�  (KK K euj\  h3j]  ]r�  j_  ]r�  ubJ��8h)�r�  }r�  (h	J��8h
X   Баженаr�  hNh]r�  (]r�  ]r�  (X   аэропОртыr�  X
   бАнтыr�  X   бОродуr�  X   бухгАлтеровr�  X   вероисповЕданиеr�  X   граждАнствоr�  X
   дефИсr�  X   диспансЕрr�  X   договорЁнностьr�  X   докумЕнтr�  X
   досУгr�  X   еретИкr�  X   жалюзИr�  X   знАчимостьr�  X   Иксыr�  X   каталОгr�  X   монолОгr�  X   квартАлr�  X   киломЕтрr�  X   кОнусыr�  X   корЫстьr�  X
   крАныr�  X   кремЕньr�  X   лЕкторыr�  X
   лыжнЯr�  X   мЕстностейr�  X   мусоропровОдr�  X   намЕрениеr�  X   нарОстr�  X   нЕдругr�  X
   недУгr�  X   некролОгr�  X   нЕнавистьr�  X   нОвостиr�  X   нОготьr�  X   Отрочествоr�  X   партЕрr�  X   портфЕльr�  X   пОручниr�  X   придАноеr�  X   призЫвr�  X
   отзЫвr�  X   свЁклаr�  X   сирОтыr�  X   срЕдстваr�  X
   созЫвr�  X   стАтуяr�  X   столЯрr�  X   тамОжняr�  X
   тОртыr�  X   цемЕнтr�  X   цЕнтнерr�  X   цепОчкаr�  X
   шАрфыr�  X
   шофЁрr�  X   экспЕртr�  X
   вернАr�  X   красИвееr�  X   красИвейшийr�  X   кУхонныйr 	  X
   ловкАr	  X   оптОвыйr	  X   прозорлИваr	  X   рядУr	  X   болтлИваr	  X   слИвовыйr	  X   брАтьсяr	  X   бралАсьr	  X
   взятьr		  X
   взялАr
	  X   взЯтьсяr	  X   взялАсьr	  X   включИтьr	  X   включИшьr	  X   включИтr	  X   включИмr	  X   влИтьсяr	  X   влилАсьr	  X   ворвАтьсяr	  X   ворвалАсьr	  X   воспринЯтьr	  X   воспринялАr	  X   воссоздАтьr	  X   воссоздалАr	  X   вручИтьr	  X   вручИтr	  X
   гнАтьr	  X
   гналАr	  X   гнАтьсяr	  X   гналАсьr	  X   добрАтьr	  X   добралАr 	  X   добрАтьсяr!	  X   добралАсьr"	  X   дождАтьсяr#	  X   дождалАсьr$	  X   дозвонИтьсяr%	  X   дозвонИтсяr&	  X   дозвонЯтсяr'	  X   дозИроватьr(	  X
   ждатьr)	  X
   ждалАr*	  X   жИтьсяr+	  X   жилОсьr,	  X   закУпоритьr-	  X   занЯтьr.	  X
   зАнялr/	  X   занялАr0	  X   зАнялоr1	  X   зАнялиr2	  X   заперЕтьr3	  X   заперлАr4	  X   заперЕтьсяr5	  X   заперлАсьr6	  X
   зватьr7	  X
   звалАr8	  X   звонИтьr9	  X   звонИшьr:	  X   звонИтr;	  X   звонИмr<	  X   исчЕрпатьr=	  X   клАстьr>	  X
   клАлаr?	  X   клЕитьr@	  X   крАстьсяrA	  X   крАласьrB	  X
   лгатьrC	  X
   лгалАrD	  X   литьrE	  X   лилАrF	  X   лИтьсяrG	  X   лилАсьrH	  X   наврАтьrI	  X   навралАrJ	  X   наделИтьrK	  X   наделИтrL	  X   надорвАтьсяrM	  X   надорвалАсьrN	  X   назвАтьсяrO	  X   назвалАсьrP	  X   накренИтьсяrQ	  X   накренИтсяrR	  X   налИтьrS	  X   налилАrT	  X   нарвАтьrU	  X   нарвалАrV	  X   насорИтьrW	  X   насорИтrX	  X   начАтьrY	  X
   нАчалrZ	  X   началАr[	  X   нАчалиr\	  X   обзвонИтьr]	  X   обзвонИтr^	  X   облегчИтьr_	  X   облегчИтr`	  X   облИтьсяra	  X   облилАсьrb	  X   обнЯтьсяrc	  X   обнялАсьrd	  X   обогнАтьre	  X   обогналАrf	  X   ободрАтьrg	  X   ободралАrh	  X   ободрИтьri	  X   ободрИтьсяrj	  X   ободрИшьсяrk	  X   обострИтьrl	  X   одолжИтьrm	  X   одолжИтrn	  X   озлОбитьro	  X   оклЕитьrp	  X   окружИтьrq	  X   окружИтrr	  X   опломбировАтьrs	  X   формировАтьrt	  X   нормировАтьru	  X   сортировАтьrv	  X   премировАтьrw	  X   опОшлитьrx	  X   освЕдомитьсяry	  X   освЕдомишьсяrz	  X   отбЫтьr{	  X   отбылАr|	  X   отдАтьr}	  X   отдалАr~	  X   откУпоритьr	  X   откУпорилr�	  X   отозвАтьr�	  X   отозвалАr�	  X   отозвАтьсяr�	  X   отозвалАсьr�	  X   перезвонИтьr�	  X   перезвонИтr�	  X   перелИтьr�	  X   перелилАr�	  X   плодоносИтьr�	  X   повторИтьr�	  X   повторИтr�	  X   позвАтьr�	  X   позвалАr�	  X   позвонИтьr�	  X   позвонИшьr�	  X   позвонИтr�	  X   полИтьr�	  X   полилАr�	  X   положИтьr�	  X   положИлr�	  X   понЯтьr�	  X   понялАr�	  X   послАтьr�	  X   послАлаr�	  X   прибЫтьr�	  X   прИбылr�	  X   прибылАr�	  X   прИбылоr�	  X   принЯтьr�	  X   прИнялr�	  X   прИнялиr�	  X   принялАr�	  X   принУдитьr�	  X
   рвАтьr�	  X
   рвалАr�	  X   сверлИтьr�	  X   сверлИшьr�	  X   сверлИтr�	  X
   снЯтьr�	  X
   снялАr�	  X   создАтьr�	  X   создалАr�	  X   сорвАтьr�	  X   сорвалАr�	  X   сорИтьr�	  X
   сорИтr�	  X   убрАтьr�	  X   убралАr�	  X   убыстрИтьr�	  X   углубИтьr�	  X   укрепИтьr�	  X   укрепИтr�	  X   чЕрпатьr�	  X   щемИтьr�	  X
   щемИтr�	  X   щЁлкатьr�	  X   балОванныйr�	  X   включЁнныйr�	  X   включЁнr�	  X   низведЁнныйr�	  X   довезЁнныйr�	  X   зАгнутыйr�	  X   зАнятыйr�	  X   занятАr�	  X   зАпертыйr�	  X   запертАr�	  X   заселЁнныйr�	  X   заселенАr�	  X   избалОванныйr�	  X   балОванныйr�	  X   кормЯщийr�	  X   кровоточАщийr�	  X   молЯщийr�	  X   нажИвшийr�	  X   нАжитыйr�	  X   нажитАr�	  X   налИвшийr�	  X   налитАr�	  X   нанЯвшийся	r�	  X   начАвшийr�	  X   нАчатыйr�	  X   низведЁнныйr�	  X   низведЁнr�	  X   включЁнныйr�	  X   ободрЁнныйr�	  X   ободрЁнr�	  X   ободренАr�	  X   обострЁнныйr�	  X   отключЁнныйr�	  X   определЁнныйr�	  X   определЁнr�	  X   отключЁнныйr�	  X   повторЁнныйr�	  X   поделЁнныйr�	  X   понЯвшийr�	  X   прИнятыйr�	  X   приручЁнныйr�	  X   прожИвшийr�	  X   снЯтыйr�	  X
   снятАr�	  X   сОгнутыйr�	  X   балУясьr�	  X   закУпоривr�	  X
   начАвr�	  X   начАвшисьr�	  X
   отдАвr�	  X   поднЯвr�	  X
   понЯвr�	  X   прибЫвr�	  X   вОвремяr�	  X   добелАr�	  X   дОверхуr�	  X   донЕльзяr�	  X   дОнизуr�	  X   дОсухаr�	  X   завИдноr�	  X   зАгодяr�	  X   зАсветлоr�	  X   зАтемноr�	  X   красИвееr�	  X   навЕрхr�	  X   надОлгоr�	  X   ненадОлгоr�	  e]r�	  ej?  }r�	  (j�	  ]r�	  (KK K ej�  ]r�	  (KK Kej	  ]r 
  (KK K ej�	  ]r
  (KK K ejT	  ]r
  (KK K ej	  ]r
  (KKKej�	  ]r
  (KK K ej�	  ]r
  (KK Kej#	  ]r
  (KK K ej{	  ]r
  (KK K ejX	  ]r
  (KK K ej�	  ]r	
  (K KKej�	  ]r

  (KK K ej�  ]r
  (KK Kej�	  ]r
  (KK K ej�  ]r
  (K KKejW	  ]r
  (KK K ejN	  ]r
  (KK K ej�	  ]r
  (KK Kej*	  ]r
  (KK K ej�  ]r
  (K KKej�  ]r
  (KK Kej�	  ]r
  (KK Kej�	  ]r
  (K KKejU	  ]r
  (KK K euj\  j8	  j]  ]r
  j_  ]r
  ubJ��h)�r
  }r
  (h	J��h
X   Sergei.r
  hNh]r
  (]r
  ]r
  (j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j 	  j	  j	  j	  j	  j	  j	  j	  j	  j		  j
	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j 	  j!	  j"	  j#	  j$	  j%	  j&	  j'	  j(	  j)	  j*	  j+	  j,	  j-	  j.	  j/	  j0	  j1	  j2	  j3	  j4	  j5	  j6	  j7	  j8	  j9	  j:	  j;	  j<	  j=	  j>	  j?	  j@	  jA	  jB	  jC	  jD	  jE	  jF	  jG	  jH	  jI	  jJ	  jK	  jL	  jM	  jN	  jO	  jP	  jQ	  jR	  jS	  jT	  jU	  jV	  jW	  jX	  jY	  jZ	  j[	  j\	  j]	  j^	  j_	  j`	  ja	  jb	  jc	  jd	  je	  jf	  jg	  jh	  ji	  jj	  jk	  jl	  jm	  jn	  jo	  jp	  jq	  jr	  js	  jt	  ju	  jv	  jw	  jx	  jy	  jz	  j{	  j|	  j}	  j~	  j	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  e]r
  ej?  }r 
  j\  j�	  j]  ]r!
  j_  ]r"
  ubJ�o�h)�r#
  }r$
  (h	J�o�h
X   Миша Репинr%
  hNh]r&
  (]r'
  ]r(
  (j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j 	  j	  j	  j	  j	  j	  j	  j	  j	  j		  j
	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j 	  j!	  j"	  j#	  j$	  j%	  j&	  j'	  j(	  j)	  j*	  j+	  j,	  j-	  j.	  j/	  j0	  j1	  j2	  j3	  j4	  j5	  j6	  j7	  j8	  j9	  j:	  j;	  j<	  j=	  j>	  j?	  j@	  jA	  jB	  jC	  jD	  jE	  jF	  jG	  jH	  jI	  jJ	  jK	  jL	  jM	  jN	  jO	  jP	  jQ	  jR	  jS	  jT	  jU	  jV	  jW	  jX	  jY	  jZ	  j[	  j\	  j]	  j^	  j_	  j`	  ja	  jb	  jc	  jd	  je	  jf	  jg	  jh	  ji	  jj	  jk	  jl	  jm	  jn	  jo	  jp	  jq	  jr	  js	  jt	  ju	  jv	  jw	  jx	  jy	  jz	  j{	  j|	  j}	  j~	  j	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  e]r)
  ej?  }r*
  (j'	  ]r+
  (KK K ej�	  ]r,
  (KK K ejB	  ]r-
  (K KKej�  ]r.
  (KK K ej�	  ]r/
  (KK K ej�	  ]r0
  (KK K ej�  ]r1
  (KK K ej	  ]r2
  (KK Kej�	  ]r3
  (KK K ejg	  ]r4
  (KK K ej�  ]r5
  (KK K ej�	  ]r6
  (KK K ej�	  ]r7
  (KK Kej�  ]r8
  (KK K ej�	  ]r9
  (KK K ej�	  ]r:
  (KK Kej�	  ]r;
  (KK K ejq	  ]r<
  (KK K ej�	  ]r=
  (K KKej�	  ]r>
  (KK K ej�  ]r?
  (KK K ej�  ]r@
  (KK K ej�  ]rA
  (KK K ej?	  ]rB
  (KK Kej�	  ]rC
  (KK Kej	  ]rD
  (KK KejX	  ]rE
  (KK KejG	  ]rF
  (KK K ej6	  ]rG
  (KK K ej�  ]rH
  (KK K ej�  ]rI
  (KK K ej�	  ]rJ
  (KK K ej�	  ]rK
  (KK K ejR	  ]rL
  (K KKej�	  ]rM
  (KK Kej	  ]rN
  (KK K ej�  ]rO
  (KK K ej�	  ]rP
  (KK K ej�  ]rQ
  (KK K ej�  ]rR
  (KK K ej�	  ]rS
  (KK K ej4	  ]rT
  (KK K ej�	  ]rU
  (KK K ej+	  ]rV
  (KK K ejx	  ]rW
  (KK K ej	  ]rX
  (KK Keuj\  j�	  j]  ]rY
  j_  ]rZ
  ubJ��"6h)�r[
  }r\
  (h	J��"6h
X   Rafatdinr]
  hNh]r^
  (]r_
  ]r`
  (j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j 	  j	  j	  j	  j	  j	  j	  j	  j	  j		  j
	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j	  j 	  j!	  j"	  j#	  j$	  j%	  j&	  j'	  j(	  j)	  j*	  j+	  j,	  j-	  j.	  j/	  j0	  j1	  j2	  j3	  j4	  j5	  j6	  j7	  j8	  j9	  j:	  j;	  j<	  j=	  j>	  j?	  j@	  jA	  jB	  jC	  jD	  jE	  jF	  jG	  jH	  jI	  jJ	  jK	  jL	  jM	  jN	  jO	  jP	  jQ	  jR	  jS	  jT	  jU	  jV	  jW	  jX	  jY	  jZ	  j[	  j\	  j]	  j^	  j_	  j`	  ja	  jb	  jc	  jd	  je	  jf	  jg	  jh	  ji	  jj	  jk	  jl	  jm	  jn	  jo	  jp	  jq	  jr	  js	  jt	  ju	  jv	  jw	  jx	  jy	  jz	  j{	  j|	  j}	  j~	  j	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  j�	  e]ra
  ej?  }rb
  (j�	  ]rc
  (K KKejc	  ]rd
  (KK K ej�	  ]re
  (KK K euj\  j�  j]  ]rf
  j�	  aj_  ]rg
  ubJK��h)�rh
  }ri
  (h	JK��h
X   Philipprj
  hNh]rk
  (]rl
  ]rm
  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rn
  ej?  }ro
  (j  ]rp
  (KK K ej;  ]rq
  (KKKej�  ]rr
  (KK K ejJ  ]rs
  (K KKejH  ]rt
  (KK Kej�  ]ru
  (KK K ej�  ]rv
  (KK K ej�  ]rw
  (K KKeje  ]rx
  (K KK ej�  ]ry
  (KK K ej�  ]rz
  (K KKej�  ]r{
  (KK K ejp  ]r|
  (KK K ejr  ]r}
  (KK K ej  ]r~
  (KK K ej@  ]r
  (KK K ejy  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (K KKejX  ]r�
  (KK Kej  ]r�
  (KK K ej�  ]r�
  (KK K ejD  ]r�
  (KK K ej�  ]r�
  (KK K ejs  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (K KK ej  ]r�
  (KK K ej�  ]r�
  (KK K euj\  j�  j]  ]r�
  j_  ]r�
  j�  aubJ%��h)�r�
  }r�
  (h	J%��h
X   Susannar�
  hNh]r�
  (]r�
  ]r�
  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  j{  j|  e]r�
  ej?  }r�
  (ji  ]r�
  (KK K ejK  ]r�
  (KK K ejV  ]r�
  (KK K ejD  ]r�
  (KK K ej  ]r�
  (KK K ejw  ]r�
  (KK K ej�  ]r�
  (KK K ej<  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej-  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK Kej�  ]r�
  (KK K eja  ]r�
  (KK K ej�  ]r�
  (KK K ejd  ]r�
  (KK K ejq  ]r�
  (KK K ej�  ]r�
  (KK K ej=  ]r�
  (KK K ejG  ]r�
  (KK K ejN  ]r�
  (KK K ej�  ]r�
  (KK K ejR  ]r�
  (KK K ej�  ]r�
  (KK Kej  ]r�
  (KK K ej  ]r�
  (KK K ej�  ]r�
  (KK K ejb  ]r�
  (KK K ejx  ]r�
  (KK K ej2  ]r�
  (KK Kejd  ]r�
  (KK K ej�  ]r�
  (KK K ej~  ]r�
  (KK K ejU  ]r�
  (KK K ej�  ]r�
  (KK K eju  ]r�
  (KK Kej�  ]r�
  (KK K ej]  ]r�
  (KK K ej�  ]r�
  (KK K ej,  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ejY  ]r�
  (KK K ej�  ]r�
  (KK K ej  ]r�
  (KK K ej  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ejo  ]r�
  (KK K ej�  ]r�
  (KK K ej
  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ejZ  ]r�
  (KK K ejz  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej  ]r�
  (KK K ej^  ]r�
  (KK K ej�  ]r�
  (KK K ejw  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ejp  ]r�
  (KK K ej�  ]r�
  (KK KejI  ]r�
  (KK K ej�  ]r�
  (KK K ejl  ]r�
  (KK K euj\  jw  j]  ]r�
  (j<  j�  j2  ju  ej_  ]r�
  (j�  j�  j�  j�  j�  j  j  j�  j�  j,  j�  j�  j  j  j�  j�  j�  jZ  jz  j�  j�  jw  eubJע~h)�r�
  }r�
  (h	Jע~h
X   Vitaliyr�
  hNh]r�
  (]r�
  ]r�
  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�
  ej?  }r�
  j\  j3  j]  ]r�
  j_  ]r�
  ubJ�n�h)�r�
  }r�
  (h	J�n�h
X   NoNaler�
  hNh]r�
  (]r�
  ]r�
  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�
  ej?  }r�
  (ja  ]r�
  (KK K eje  ]r�
  (KK K ejy  ]r�
  (KK K eja  ]r�
  (KK K ej�  ]r�
  (KK K ejx  ]r�
  (KK K ej�  ]r�
  (KK K ej  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r�
  (KK K ej�  ]r   (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ejw  ]r  (KK K ejn  ]r  (KK K ejd  ]r  (KK K ej!  ]r  (KK K ejx  ]r  (KK K ej�  ]r	  (KK K ej[  ]r
  (KK K ej@  ]r  (KK K ej�  ]r  (KK K ejE  ]r  (KK K ej�  ]r  (KK K ej"  ]r  (KK K ej  ]r  (KK K ej  ]r  (KK K ejM  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K eju  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej  ]r  (KK K ej  ]r  (KK K ejv  ]r  (KK K ej]  ]r  (KK K ejB  ]r  (KK K ejT  ]r  (KK K ej#  ]r   (KK K ej�  ]r!  (KK K ej|  ]r"  (KK K ej�  ]r#  (KK K ejc  ]r$  (KK K ejI  ]r%  (KK K ej
  ]r&  (KK K ej�  ]r'  (KK K ej�  ]r(  (KK K ej�  ]r)  (KK K ej]  ]r*  (KK K ej*  ]r+  (KK K ejV  ]r,  (KK K ej�  ]r-  (KK K ej  ]r.  (KK K ej�  ]r/  (KK K ej�  ]r0  (KK K ej  ]r1  (KK K ej�  ]r2  (KK K ej�  ]r3  (KK K ejR  ]r4  (KK K ejn  ]r5  (KK K ej�  ]r6  (KK K ejz  ]r7  (KK K ej�  ]r8  (KK K ej&  ]r9  (KK K ej}  ]r:  (KK K ejG  ]r;  (KK K ej�  ]r<  (KK K ej�  ]r=  (KK K ejT  ]r>  (KK K ejz  ]r?  (KK K ej4  ]r@  (KK K ejt  ]rA  (KK K ej�  ]rB  (KK K ejX  ]rC  (KK K ej�  ]rD  (KK K ejZ  ]rE  (KK K ej�  ]rF  (KK K euj\  j  j]  ]rG  ja  aj_  ]rH  ubJ���/h)�rI  }rJ  (h	J���/h
X   ▪️rK  hNh]rL  (]rM  ]rN  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rO  ej?  }rP  jZ  ]rQ  (KK K esj\  jL  j]  ]rR  j_  ]rS  ubJ\�!h)�rT  }rU  (h	J\�!h
X   donny3zMrV  hNh]rW  (]rX  ]rY  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rZ  ej?  }r[  (je  ]r\  (KK K ej@  ]r]  (KK K euj\  j;  j]  ]r^  jG  aj_  ]r_  (jA  je  j@  eubJs`Gh)�r`  }ra  (h	Js`Gh
X   Margorb  hNh]rc  (]rd  ]re  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rf  ej?  }rg  (j�  ]rh  (KK Kej  ]ri  (KK Kej�  ]rj  (KK K ejY  ]rk  (KK Kej�  ]rl  (KK Keuj\  jJ  j]  ]rm  j  aj_  ]rn  ubJ1�3h)�ro  }rp  (h	J1�3h
X   Евгенияrq  hNh]rr  (]rs  ]rt  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]ru  ej?  }rv  j\  jA  j]  ]rw  j_  ]rx  ubJnQ�h)�ry  }rz  (h	JnQ�h
X   Dashar{  hNh]r|  (]r}  ]r~  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r  ej?  }r�  (j�  ]r�  (KK K ej�  ]r�  (KK K eje  ]r�  (KK K ejx  ]r�  (KK K ejT  ]r�  (KK K ej�  ]r�  (KK K ej_  ]r�  (KK K ej	  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej[  ]r�  (KK K ejY  ]r�  (KK K ejV  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej   ]r�  (KK K ej�  ]r�  (K KKej�  ]r�  (KK K ej�  ]r�  (KK K ejU  ]r�  (KK K ej�  ]r�  (KK K ejI  ]r�  (KK K ej  ]r�  (KK K ejR  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejQ  ]r�  (KK K ejd  ]r�  (KK K ej�  ]r�  (K KKej(  ]r�  (KK K ej�  ]r�  (K KKejK  ]r�  (K KKej�  ]r�  (KK K ejP  ]r�  (KK K ejt  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej  ]r�  (KK K euj\  j�  j]  ]r�  j�  aj_  ]r�  ubJp�,9h)�r�  }r�  (h	Jp�,9h
X   Annr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (jZ  ]r�  (KK Kej�  ]r�  (KKK ejq  ]r�  (KK K ej[  ]r�  (KK Kej'  ]r�  (KK K ej�  ]r�  (KKKej�  ]r�  (KK K ej4  ]r�  (KK K ej�  ]r�  (KK K ejq  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ejn  ]r�  (KK K ejQ  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej{  ]r�  (KK K ejs  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej
  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ejx  ]r�  (KK K ejB  ]r�  (KK Kej�  ]r�  (KK Kej)  ]r�  (KK K ejM  ]r�  (KK K ejw  ]r�  (KK K ej�  ]r�  (KK K ej_  ]r�  (KK K ejX  ]r�  (KK K ej�  ]r�  (KK K ejm  ]r�  (KK Keju  ]r�  (KK K ej  ]r�  (KK KejC  ]r�  (KK K ej  ]r�  (KK K ejY  ]r�  (KK K ej*  ]r�  (KK K ej\  ]r�  (KK K ej[  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ejf  ]r�  (KK Kej�  ]r�  (KK K ejx  ]r�  (KK Kej�  ]r�  (KK K ejT  ]r�  (KK Kej}  ]r�  (KK K ejN  ]r�  (KK Kej  ]r�  (KK K ejJ  ]r�  (KK Kej�  ]r�  (KK Kej  ]r�  (KK Kej`  ]r�  (KK K ej�  ]r�  (KK K ej9  ]r�  (KK Kej�  ]r�  (KK K ej|  ]r�  (KK Kej�  ]r�  (KK K ej-  ]r�  (KK K ej,  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ejN  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK Kejk  ]r�  (KK K ejd  ]r�  (KK K ej�  ]r�  (KK K ejF  ]r�  (KK K ej  ]r�  (KK K ej;  ]r�  (KK Kej�  ]r�  (KK K ej!  ]r   (KK K ej  ]r  (KK K ejR  ]r  (KK Kej�  ]r  (KK K ej0  ]r  (KK K eje  ]r  (KK Kej�  ]r  (KK K ej  ]r  (KK K ejh  ]r  (KK Kejr  ]r	  (KK K ej�  ]r
  (KK K ejj  ]r  (KK K ej  ]r  (KK K ejI  ]r  (KK Kej  ]r  (KK K ej^  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ejh  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej/  ]r  (KK K euj\  j�  j]  ]r  (jJ  j�  ej_  ]r  (j�  jN  eubJ�,h)�r  }r  (h	J�,h
X
   Ксюшаr  hNh]r  (]r   ]r!  (jG  jH  jI  jJ  jK  jL  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jZ  j[  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r"  ej?  }r#  (j  ]r$  (KK Kej`  ]r%  (KK K ej�  ]r&  (KK K ejK  ]r'  (KKKej�  ]r(  (KK K ejU  ]r)  (KK K ej�  ]r*  (KKK ej  ]r+  (KK K ej�  ]r,  (KK K ejh  ]r-  (KK K ejt  ]r.  (KK K ej�  ]r/  (KK K ej�  ]r0  (KK K ej  ]r1  (KK K ej  ]r2  (KK Kej  ]r3  (KK K ejs  ]r4  (KK K ejv  ]r5  (KK Kej  ]r6  (KK K ej  ]r7  (KK K ej  ]r8  (KK K ej�  ]r9  (KK Kej�  ]r:  (KKKej\  ]r;  (KK K ej  ]r<  (KK K ejg  ]r=  (KK K ej�  ]r>  (KK K ejJ  ]r?  (KKKej
  ]r@  (KK K ej^  ]rA  (KK K ejX  ]rB  (KK K ej�  ]rC  (K KKej�  ]rD  (K KKej[  ]rE  (KK Kejz  ]rF  (KK K ej�  ]rG  (KK K ejQ  ]rH  (KK K ej0  ]rI  (KK K ejZ  ]rJ  (KKK ej{  ]rK  (KK K ejM  ]rL  (KK K ej   ]rM  (KK K ejr  ]rN  (KK K ejI  ]rO  (KK K ejx  ]rP  (KK K ej   ]rQ  (KK K ej  ]rR  (KK K ej�  ]rS  (K KKejV  ]rT  (KK K ej�  ]rU  (KK K ej-  ]rV  (KK K ej�  ]rW  (KK Kej�  ]rX  (KK Kejr  ]rY  (KK K ej�  ]rZ  (KK K ej�  ]r[  (KK K ej  ]r\  (KK K ejL  ]r]  (KK K ejI  ]r^  (KK Kej7  ]r_  (KK K ej  ]r`  (KK K ejN  ]ra  (KK Kej+  ]rb  (KK K ej�  ]rc  (KK Kej�  ]rd  (KK Kej=  ]re  (KK K ejk  ]rf  (KK K ej�  ]rg  (KK K ej!  ]rh  (KK K ej�  ]ri  (KK K ej%  ]rj  (KK K ej�  ]rk  (KK K ej�  ]rl  (KK K ej�  ]rm  (K KKej�  ]rn  (KK K ejT  ]ro  (KK K ej�  ]rp  (K KKejt  ]rq  (KK Kej�  ]rr  (KK K ej  ]rs  (KK K ej�  ]rt  (KK Kejn  ]ru  (KK K ej4  ]rv  (KK K ej�  ]rw  (KK K ej�  ]rx  (KK K ejW  ]ry  (KK K ejc  ]rz  (KK K ejS  ]r{  (KK KejF  ]r|  (KK Kejm  ]r}  (KK K ej  ]r~  (KK Kej�  ]r  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej*  ]r�  (KK K ejH  ]r�  (KK KejU  ]r�  (KK Kej  ]r�  (KK K ejA  ]r�  (KK Keja  ]r�  (KK Kej	  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK K ej/  ]r�  (K KKej�  ]r�  (KK K ejv  ]r�  (KK K ej@  ]r�  (KK K ej�  ]r�  (KK Kejx  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK Kej_  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ejj  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK Kej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejc  ]r�  (KK K ejd  ]r�  (KK K ejW  ]r�  (KK K ejY  ]r�  (KK K ejb  ]r�  (KK K ejw  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejq  ]r�  (KK K euj\  j�  j]  ]r�  jT  aj_  ]r�  (j  j0  jh  jM  j  j  j  jg  j\  jY  eubJ��7h)�r�  }r�  (h	J��7h
X   еся отвалиr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (j�  ]r�  (KK K ejR  ]r�  (KK K ejX  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej5  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejd  ]r�  (KK K ej�  ]r�  (KK K ejt  ]r�  (KK K ej�  ]r�  (KK K ej+  ]r�  (KK K ejZ  ]r�  (K KK ejh  ]r�  (KK K ejr  ]r�  (KK K ej$  ]r�  (KK K ejM  ]r�  (KK K ej�  ]r�  (KK K ej^  ]r�  (KK K ej_  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejT  ]r�  (KK K ejp  ]r�  (K KKejb  ]r�  (KK K ejt  ]r�  (KK K ej�  ]r�  (KK K eju  ]r�  (K KKej�  ]r�  (KK K ejH  ]r�  (KK K ej  ]r�  (KK K ej6  ]r�  (KK K ej
  ]r�  (KK K ej.  ]r�  (KK K ej"  ]r�  (KK K ejV  ]r�  (KK K ej�  ]r�  (KK K ejs  ]r�  (KK K ej8  ]r�  (KK K ejU  ]r�  (K KKejc  ]r�  (KK K ejy  ]r�  (KK K ej�  ]r�  (KK K ejz  ]r�  (KK K ej}  ]r�  (KK K ejg  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ejs  ]r�  (K KKej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej\  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K euj\  jy  j]  ]r�  j_  ]r�  ubJHK�h)�r�  }r�  (h	JHK�h
X
   Deathstorer�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (j\  ]r�  (KK K ej?  ]r�  (K KKejR  ]r�  (KK KejS  ]r�  (KK K ej  ]r�  (KK Kej�  ]r�  (KK K ejO  ]r�  (KK K ejY  ]r   (KK Kej|  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK Kejl  ]r  (KK K ejq  ]r  (KK Keuj\  j�  j]  ]r  j_  ]r  ubJӚmh)�r  }r	  (h	JӚmh
X   owlr
  hNh]r  (]r  ]r  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r  ej?  }r  j\  jg  j]  ]r  j_  ]r  ubJ
ߝh)�r  }r  (h	J
ߝh
X   Матвейr  hNh]r  (]r  ]r  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r  ej?  }r  j\  j`  j]  ]r  j_  ]r  ubJ4�l.h)�r  }r  (h	J4�l.h
X   ЫЫЫЫЫЫЫr  hNh]r  (]r   ]r!  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r"  ej?  }r#  j�  ]r$  (KK K esj\  j�  j]  ]r%  j_  ]r&  ubJ�x�2h)�r'  }r(  (h	J�x�2h
X   dat girlr)  hNh]r*  (]r+  ]r,  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r-  ej?  }r.  j\  jn  j]  ]r/  jn  aj_  ]r0  ubJ��/h)�r1  }r2  (h	J��/h
X   Dianar3  hNh]r4  (]r5  ]r6  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r7  ej?  }r8  (jz  ]r9  (KK K ej8  ]r:  (K KKej  ]r;  (KK K ej�  ]r<  (KK K ej�  ]r=  (KK Kejz  ]r>  (KK Keuj\  j�  j]  ]r?  j�  aj_  ]r@  j�  aubJ���h)�rA  }rB  (h	J���h
X   jjrC  hNh]rD  (]rE  ]rF  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rG  ej?  }rH  j\  j�  j]  ]rI  j_  ]rJ  ubJ�8� h)�rK  }rL  (h	J�8� h
X   RennrM  hNh]rN  (]rO  ]rP  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rQ  ej?  }rR  (j�  ]rS  (KK K ej�  ]rT  (KK Keuj\  j  j]  ]rU  j  aj_  ]rV  j�  aubJC(�=h)�rW  }rX  (h	JC(�=h
X4   𝙲𝚒𝚝𝚘𝚏𝚝𝚑𝚎𝚆𝚆 ( 𝙴*** )rY  hNh]rZ  (]r[  ]r\  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r]  ej?  }r^  (jW  ]r_  (KK Kej�  ]r`  (KK K euj\  j�  j]  ]ra  j�  aj_  ]rb  jW  aubJO=4;h)�rc  }rd  (h	JO=4;h
X   Julyre  hNh]rf  (]rg  ]rh  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]ri  ej?  }rj  (jH  ]rk  (KK K ej]  ]rl  (KK K ejY  ]rm  (KK K ej=  ]rn  (KK K eje  ]ro  (KK K ej�  ]rp  (KK K ej�  ]rq  (KK K ej�  ]rr  (KK K ejU  ]rs  (KK K eja  ]rt  (KK K eji  ]ru  (KK K ej/  ]rv  (KK K ej�  ]rw  (KK K ej�  ]rx  (KK K ej�  ]ry  (KK K euj\  jt  j]  ]rz  j_  ]r{  ubJ>�lh)�r|  }r}  (h	J>�lh
X
   Алинаr~  hNh]r  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  j�  ]r�  (KK K esj\  j{  j]  ]r�  j_  ]r�  ubJ�k�Ch)�r�  }r�  (h	J�k�Ch
X   Выжатый помидорr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  j\  j�  j]  ]r�  j_  ]r�  ubJ*6�3h)�r�  }r�  (h	J*6�3h
X   твой кавалерr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (j�  ]r�  (KK K ej]  ]r�  (KK Kejh  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej;  ]r�  (KK K ej9  ]r�  (KK K ej�  ]r�  (KK K ejS  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejw  ]r�  (KK K ejn  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejc  ]r�  (KK K ejP  ]r�  (KK Kej+  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK Kej@  ]r�  (KK Kej�  ]r�  (KK KejQ  ]r�  (KK KejC  ]r�  (KK Kej�  ]r�  (KK Keje  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK Kej  ]r�  (KK K ejV  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ejb  ]r�  (KK K ej�  ]r�  (KK K ejL  ]r�  (KK K ej2  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejK  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (K KK ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejg  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejS  ]r�  (KK K ej�  ]r�  (KK K ejU  ]r�  (KK K ej,  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejI  ]r�  (KK K euj\  j�  j]  ]r�  j�  aj_  ]r�  ubJJ�h)�r�  }r�  (h	JJ�h
X   Ленаr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  j\  jk  j]  ]r�  j_  ]r�  ubJ@f[Ch)�r�  }r�  (h	J@f[Ch
X
   suzy❣️r�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  j\  jF  j]  ]r�  j_  ]r�  ubJ�\'h)�r�  }r�  (h	J�\'h
X	   Ekaterinar�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (jy  ]r�  (KK K ejH  ]r�  (KK Kejh  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ej'  ]r�  (KK Kej  ]r�  (KK K ej  ]r�  (KK K ej#  ]r�  (KK K ej&  ]r�  (KK Kej�  ]r   (KK K eji  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K eju  ]r  (KK K ej  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej%  ]r  (KK K euj\  jA  j]  ]r	  j_  ]r
  j#  aubJ���h)�r  }r  (h	J���h
X   Йоr  hNh]r  (]r  ]r  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r  ej?  }r  (jz  ]r  (KK K ej?  ]r  (KK Kej�  ]r  (KK K ej'  ]r  (KK Kej  ]r  (KK K ej]  ]r  (KK Kejd  ]r  (KK K ej�  ]r  (KK K euj\  j�  j]  ]r  jz  aj_  ]r  j�  aubJ�Y&6h)�r  }r  (h	J�Y&6h
X   Veronikar  hNh]r   (]r!  ]r"  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r#  ej?  }r$  (j�  ]r%  (KK KejL  ]r&  (K KKej�  ]r'  (KK Kej�  ]r(  (KK Kej  ]r)  (KK Keuj\  jY  j]  ]r*  (j�  jY  ej_  ]r+  j�  aubJS1.h)�r,  }r-  (h	JS1.h
X   Valeriar.  hNh]r/  (]r0  ]r1  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r2  ej?  }r3  (je  ]r4  (KK K eji  ]r5  (KK K ej�  ]r6  (KK K ejP  ]r7  (KK Kejo  ]r8  (KK K ej�  ]r9  (KK K ej  ]r:  (KK K ejU  ]r;  (KK K ejU  ]r<  (KK K ejI  ]r=  (KK K ej�  ]r>  (KK K ej  ]r?  (KK K ej2  ]r@  (KK Kej  ]rA  (KK K ejf  ]rB  (KK K ej�  ]rC  (KK K ej^  ]rD  (KK K ej�  ]rE  (KK K ej  ]rF  (KK K ejC  ]rG  (KK K ej�  ]rH  (KK K ej?  ]rI  (KK K ejN  ]rJ  (KK K ej�  ]rK  (KK K ej`  ]rL  (KK K ejv  ]rM  (KK K ej   ]rN  (KK K ej  ]rO  (KK K ej%  ]rP  (KK K ej  ]rQ  (KK K ejV  ]rR  (KK K eja  ]rS  (KK K ej�  ]rT  (KK K ej  ]rU  (KK Kej�  ]rV  (KK K ejs  ]rW  (KK K ej^  ]rX  (KK K ejp  ]rY  (KK K ej  ]rZ  (KK K ejO  ]r[  (KK K ejl  ]r\  (KK K ejz  ]r]  (KK K ejj  ]r^  (KK K ej�  ]r_  (KK K ej�  ]r`  (KK K ejR  ]ra  (KK Kej7  ]rb  (KK K ej�  ]rc  (KK K ej!  ]rd  (KK K eja  ]re  (KK Kej�  ]rf  (KK Kej�  ]rg  (KK Kej�  ]rh  (KK Keuj\  j   j]  ]ri  j_  ]rj  j�  aubJ@�aAh)�rk  }rl  (h	J@�aAh
X
   Stephendorrm  hNh]rn  (]ro  ]rp  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rq  ej?  }rr  j\  j�  j]  ]rs  j_  ]rt  ubJ��V=h)�ru  }rv  (h	J��V=h
X   Olyarw  hNh]rx  (]ry  ]rz  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r{  ej?  }r|  (j�  ]r}  (KK K ej  ]r~  (KK K ejZ  ]r  (K KKeuj\  j2  j]  ]r�  (j�  j  ej_  ]r�  jZ  aubJ[�`*h)�r�  }r�  (h	J[�`*h
X   Аидаr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  j\  j�  j]  ]r�  j_  ]r�  ubJ)V)<h)�r�  }r�  (h	J)V)<h
X   Dariar�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  j\  j.  j]  ]r�  j_  ]r�  ubJ��Sh)�r�  }r�  (h	J��Sh
X   Kasiar�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (j`  ]r�  (KK K ejK  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ejz  ]r�  (KK K ej{  ]r�  (KK K ejf  ]r�  (KK K ejd  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K eje  ]r�  (KK K ejx  ]r�  (KK K ejv  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej8  ]r�  (KK K ej=  ]r�  (KK K ej�  ]r�  (KK K ej>  ]r�  (KK K ej�  ]r�  (KK K ej|  ]r�  (KK K ej3  ]r�  (KK K ejG  ]r�  (KK K ej�  ]r�  (KK K ejW  ]r�  (KK K ej`  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej  ]r�  (KK K ejD  ]r�  (KK K ej�  ]r�  (KK K ejt  ]r�  (KK K ejV  ]r�  (KK K ej  ]r�  (KK K ej-  ]r�  (KK K ej�  ]r�  (KK K ejn  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K eju  ]r�  (KK K ej�  ]r�  (KK K ejw  ]r�  (KK K ej�  ]r�  (KK K ejJ  ]r�  (KK K ej�  ]r�  (KK Kejk  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ejG  ]r�  (KK K ej^  ]r�  (KK K ejj  ]r�  (KK K eju  ]r�  (KK K ej_  ]r�  (KK K ej�  ]r�  (KK Keja  ]r�  (KK K ej*  ]r�  (KK K ejr  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK KejT  ]r�  (KK K euj\  j�  j]  ]r�  j_  ]r�  (j�  j=  jn  j_  eubJw�7h)�r�  }r�  (h	Jw�7h
X   Dr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (jq  ]r�  (KK K ej;  ]r�  (KK Kej  ]r�  (KK K ej  ]r�  (KK K ejV  ]r�  (KK K eju  ]r�  (KK K ej�  ]r�  (KK K ejs  ]r�  (KK K ejz  ]r�  (KK K ejd  ]r�  (KK K ejo  ]r�  (KK K ej�  ]r�  (KK K ej7  ]r�  (KK K ej�  ]r�  (KK K ejf  ]r�  (KK K ejg  ]r�  (KK K ejH  ]r�  (KK K ej�  ]r   (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej>  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej�  ]r	  (KK K ej�  ]r
  (KK K ej�  ]r  (KK K ejr  ]r  (KK K eji  ]r  (KK K ejZ  ]r  (KK K ej  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej&  ]r  (KK K ej�  ]r  (KK K ej�  ]r  (KK K ej@  ]r  (KK K euj\  jo  j]  ]r  j;  aj_  ]r  ubJ�h�3h)�r  }r  (h	J�h�3h
X   Никитаr  hNh]r  (]r  ]r  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r  ej?  }r  (jx  ]r   (KK Kejs  ]r!  (KK K ej`  ]r"  (KK Kej�  ]r#  (K KK ej�  ]r$  (K KKej�  ]r%  (K KKej  ]r&  (KK K ej�  ]r'  (KK Kej  ]r(  (KKKej  ]r)  (KK Kej�  ]r*  (K KKej   ]r+  (KK Kej�  ]r,  (KK Kejk  ]r-  (KK Kejn  ]r.  (KK Keja  ]r/  (KK KejO  ]r0  (KK K ej  ]r1  (KK Keuj\  j�  j]  ]r2  (jx  j`  j�  j  jn  ja  jO  ej_  ]r3  ubJ�X�+h)�r4  }r5  (h	J�X�+h
X   Zaikar6  hNh]r7  (]r8  ]r9  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r:  ej?  }r;  j\  j�  j]  ]r<  j_  ]r=  ubJ(EM#h)�r>  }r?  (h	J(EM#h
X   Евгенийr@  hNh]rA  (]rB  ]rC  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rD  ej?  }rE  (jn  ]rF  (KK K ej�  ]rG  (KK K ej[  ]rH  (KK K ejP  ]rI  (KK Kejm  ]rJ  (KK K ej�  ]rK  (KK K ej�  ]rL  (KK K ej2  ]rM  (KK K ej�  ]rN  (KK K ejg  ]rO  (KK Kej  ]rP  (KK K ej�  ]rQ  (KK K ejO  ]rR  (KK KejI  ]rS  (KK K ej�  ]rT  (KK K ej�  ]rU  (KK K ejw  ]rV  (KK K ej�  ]rW  (KK K ej�  ]rX  (KK K ej�  ]rY  (KK K ej�  ]rZ  (KK K euj\  j`  j]  ]r[  j_  ]r\  jo  aubJ�A�,h)�r]  }r^  (h	J�A�,h
X   Мариr_  hNh]r`  (]ra  ]rb  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j|  e]rc  ej?  }rd  j{  ]re  (KK K esj\  j�  j]  ]rf  j�  aj_  ]rg  j{  aubJ��0h)�rh  }ri  (h	J��0h
X   Анастасияrj  hNh]rk  (]rl  ]rm  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rn  ej?  }ro  (jF  ]rp  (KK K ej  ]rq  (KK K ejQ  ]rr  (KK K ej�  ]rs  (KK K ej(  ]rt  (KK K ejU  ]ru  (KK K ejn  ]rv  (KK K ejb  ]rw  (KK Kejw  ]rx  (KK K ejN  ]ry  (KK K eja  ]rz  (KK K ej�  ]r{  (KK K ejK  ]r|  (KK K ej  ]r}  (KK K ej:  ]r~  (KK K ejz  ]r  (KK K ejX  ]r�  (KK K ej]  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej6  ]r�  (KK Kej  ]r�  (KK K ej8  ]r�  (KK K ejf  ]r�  (KK K ej�  ]r�  (KK Kej|  ]r�  (KK K ej�  ]r�  (KK K ejJ  ]r�  (KK K ej�  ]r�  (KK K ej*  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K ej#  ]r�  (KK K eje  ]r�  (KK K ejX  ]r�  (KK K ej�  ]r�  (KK Keji  ]r�  (KK K ej  ]r�  (KK K euj\  j_  j]  ]r�  j_  aj_  ]r�  jn  aubJ��h)�r�  }r�  (h	J��h
X   mancr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  j\  j`  j]  ]r�  j_  ]r�  ubJ��|h)�r�  }r�  (h	J��|h
X   Yaroslavr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (j�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK Kej�  ]r�  (KK Keje  ]r�  (K KKej  ]r�  (KK K ejI  ]r�  (KK K ej�  ]r�  (K KKej�  ]r�  (KK K ej�  ]r�  (K KKejT  ]r�  (KK K ejo  ]r�  (KK K ej  ]r�  (KK K ej  ]r�  (KK K ej^  ]r�  (KK K ej�  ]r�  (KK Kejh  ]r�  (KK Kej�  ]r�  (KK Kejz  ]r�  (KK K ej�  ]r�  (KK K ejq  ]r�  (K KKej`  ]r�  (KK K ej%  ]r�  (KK K eji  ]r�  (KK K ej�  ]r�  (KK K eja  ]r�  (KK K ejN  ]r�  (KK K ej  ]r�  (KK K ej]  ]r�  (KK K ej�  ]r�  (KK K ejq  ]r�  (KK K ejC  ]r�  (KK K ej<  ]r�  (KK K ejm  ]r�  (KK K ej�  ]r�  (KKK ej  ]r�  (KK Kej�  ]r�  (KK K ej�  ]r�  (K KK ej�  ]r�  (KK K ejN  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ejS  ]r�  (KK Kej�  ]r�  (K KKej�  ]r�  (KK K ejb  ]r�  (KK K ejQ  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ejc  ]r�  (KK K ej  ]r�  (KK K ej  ]r�  (KK K ej  ]r�  (KK K ej�  ]r�  (KK K ejG  ]r�  (KK K ej�  ]r�  (KK K ej  ]r�  (KK K ejF  ]r�  (KK K ejw  ]r�  (KK K ej5  ]r�  (KK K ejd  ]r�  (KK K ejp  ]r�  (K KK ejy  ]r�  (KK K ej�  ]r�  (KK K euj\  jY  j]  ]r�  j_  ]r�  ubJu%!h)�r�  }r�  (h	Ju%!h
X   Димаr�  hNh]r�  (]r�  ]r�  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r�  ej?  }r�  (j�  ]r�  (KK Kej  ]r�  (KK K euj\  j  j]  ]r�  j_  ]r�  j�  aubJӮ�$h)�r�  }r�  (h	JӮ�$h
X
   Настяr�  hNh]r   (]r  ]r  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r  ej?  }r  (jR  ]r  (KK Kej>  ]r  (KK Kej�  ]r  (KK K euj\  j�  j]  ]r  j_  ]r	  (jR  j>  eubJ�R! h)�r
  }r  (h	J�R! h
X   Adelyar  hNh]r  (]r  ]r  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r  ej?  }r  (jH  ]r  (KK K ej.  ]r  (KK K ejP  ]r  (KK K ej  ]r  (KK K ejG  ]r  (KK K ejl  ]r  (KK K ej�  ]r  (KK K ej|  ]r  (KK K ej�  ]r  (KK K ej]  ]r  (KK K ej�  ]r  (K KKej,  ]r  (KK Kej�  ]r  (K KKej�  ]r  (KK Kej�  ]r   (KK Kejh  ]r!  (KK Kej�  ]r"  (KK Kej�  ]r#  (KK Kej�  ]r$  (KK Keuj\  j�  j]  ]r%  j_  ]r&  ubJ剌&h)�r'  }r(  (h	J剌&h
X   Danr)  hNh]r*  (]r+  ]r,  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r-  ej?  }r.  (jb  ]r/  (KK K ej�  ]r0  (KK K ej�  ]r1  (KK K ej�  ]r2  (KK K ej�  ]r3  (KK K ej�  ]r4  (KK K ej�  ]r5  (KK K euj\  j�  j]  ]r6  j_  ]r7  ubJ�k?h)�r8  }r9  (h	J�k?h
X
   Еленаr:  hNh]r;  (]r<  ]r=  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r>  ej?  }r?  j\  j  j]  ]r@  j_  ]rA  ubJB�h)�rB  }rC  (h	JB�h
X
   ЭлинаrD  hNh]rE  (]rF  ]rG  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rH  ej?  }rI  (j1  ]rJ  (KK K ejS  ]rK  (KK K ej`  ]rL  (KK Keuj\  j�  j]  ]rM  (jS  j`  ej_  ]rN  ubJ��u>h)�rO  }rP  (h	J��u>h
X
   ToP_KO$MO$rQ  hNh]rR  (]rS  ]rT  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rU  ej?  }rV  jL  ]rW  (KK K esj\  jS  j]  ]rX  j_  ]rY  ubJ�+�h)�rZ  }r[  (h	J�+�h
X   Wsssar\  hNh]r]  (]r^  ]r_  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]r`  ej?  }ra  j\  jS  j]  ]rb  j_  ]rc  ubJ��C>h)�rd  }re  (h	J��C>h
X   JOKERrf  hNh]rg  (]rh  ]ri  (jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  e]rj  ej?  }rk  (j!  ]rl  (KK K ejd  ]rm  (KK Kej\  ]rn  (KK Kej  ]ro  (KK K ej\  ]rp  (KK Kej  ]rq  (KK Kej�  ]rr  (KK K ej�  ]rs  (KK KejO  ]rt  (KK Keuj\  j�  j]  ]ru  j!  aj_  ]rv  j!  aubJ0V�@h)�rw  }rx  (h	J0V�@h
X   *<Qarakesek>*ry  hNh]rz  (]r{  ]r|  (X   аэропОртыr}  X
   бАнтыr~  X   бОродуr  X   бухгАлтеровr�  X   вероисповЕданиеr�  X   граждАнствоr�  X
   дефИсr�  X   диспансЕрr�  X   договорЁнностьr�  X   докумЕнтr�  X
   досУгr�  X   еретИкr�  X   жалюзИr�  X   знАчимостьr�  X   Иксыr�  X   каталОгr�  X   монолОгr�  X   квартАлr�  X   киломЕтрr�  X   кОнусыr�  X   корЫстьr�  X
   крАныr�  X   кремЕньr�  X   лЕкторыr�  X
   лыжнЯr�  X   мЕстностейr�  X   мусоропровОдr�  X   намЕрениеr�  X   нарОстr�  X   нЕдругr�  X
   недУгr�  X   некролОгr�  X   нЕнавистьr�  X   нОвостиr�  X   нОготьr�  X   Отрочествоr�  X   партЕрr�  X   портфЕльr�  X   пОручниr�  X   придАноеr�  X   призЫвr�  X
   отзЫвr�  X   свЁклаr�  X   сирОтыr�  X   срЕдстваr�  X
   созЫвr�  X   стАтуяr�  X   столЯрr�  X   тамОжняr�  X
   тОртыr�  X   цемЕнтr�  X   цЕнтнерr�  X   цепОчкаr�  X
   шАрфыr�  X
   шофЁрr�  X   экспЕртr�  X
   вернАr�  X   красИвееr�  X   красИвейшийr�  X   кУхонныйr�  X
   ловкАr�  X   оптОвыйr�  X   прозорлИваr�  X   рядУr�  X   болтлИваr�  X   слИвовыйr�  X   брАтьсяr�  X   бралАсьr�  X
   взятьr�  X
   взялАr�  X   взЯтьсяr�  X   взялАсьr�  X   включИтьr�  X   включИшьr�  X   включИтr�  X   включИмr�  X   влИтьсяr�  X   влилАсьr�  X   ворвАтьсяr�  X   ворвалАсьr�  X   воспринЯтьr�  X   воспринялАr�  X   воссоздАтьr�  X   воссоздалАr�  X   вручИтьr�  X   вручИтr�  X
   гнАтьr�  X
   гналАr�  X   гнАтьсяr�  X   гналАсьr�  X   добрАтьr�  X   добралАr�  X   добрАтьсяr�  X   добралАсьr�  X   дождАтьсяr�  X   дождалАсьr�  X   дозвонИтьсяr�  X   дозвонИтсяr�  X   дозвонЯтсяr�  X   дозИроватьr�  X
   ждатьr�  X
   ждалАr�  X   жИтьсяr�  X   жилОсьr�  X   закУпоритьr�  X   занЯтьr�  X
   зАнялr�  X   занялАr�  X   зАнялоr�  X   зАнялиr�  X   заперЕтьr�  X   заперлАr�  X   заперЕтьсяr�  X   заперлАсьr�  X
   зватьr�  X
   звалАr�  X   звонИтьr�  X   звонИшьr�  X   звонИтr�  X   звонИмr�  X   исчЕрпатьr�  X   клАстьr�  X
   клАлаr�  X   клЕитьr�  X   крАстьсяr�  X   крАласьr�  X
   лгатьr�  X
   лгалАr�  X   литьr�  X   лилАr�  X   лилАсьr�  X   наврАтьr   X   навралАr  X   наделИтьr  X   наделИтr  X   надорвАтьсяr  X   надорвалАсьr  X   назвАтьсяr  X   назвалАсьr  X   накренИтьсяr  X   накренИтсяr	  X   налИтьr
  X   налилАr  X   нарвАтьr  X   нарвалАr  X   насорИтьr  X   насорИтr  X   начАтьr  X
   нАчалr  X   началАr  X   нАчалиr  X   обзвонИтьr  X   обзвонИтr  X   облегчИтьr  X   облегчИтr  X   облИтьсяr  X   облилАсьr  X   обнЯтьсяr  X   обнялАсьr  X   обогнАтьr  X   обогналАr  X   ободрАтьr  X   ободралАr  X   ободрИтьr   X   ободрИтьсяr!  X   ободрИшьсяr"  X   обострИтьr#  X   одолжИтьr$  X   одолжИтr%  X   озлОбитьr&  X   оклЕитьr'  X   окружИтьr(  X   окружИтr)  X   опломбировАтьr*  X   формировАтьr+  X   нормировАтьr,  X   сортировАтьr-  X   премировАтьr.  X   опОшлитьr/  X   освЕдомитьсяr0  X   освЕдомишьсяr1  X   отбЫтьr2  X   отбылАr3  X   отдАтьr4  X   отдалАr5  X   откУпоритьr6  X   откУпорилr7  X   отозвАтьr8  X   отозвалАr9  X   отозвАтьсяr:  X   отозвалАсьr;  X   перезвонИтьr<  X   перезвонИтr=  X   перелИтьr>  X   перелилАr?  X   плодоносИтьr@  X   повторИтьrA  X   повторИтrB  X   позвАтьrC  X   позвалАrD  X   позвонИтьrE  X   позвонИшьrF  X   позвонИтrG  X   полИтьrH  X   полилАrI  X   положИтьrJ  X   положИлrK  X   понЯтьrL  X   понялАrM  X   послАтьrN  X   послАлаrO  X   прибЫтьrP  X   прИбылrQ  X   прибылАrR  X   прИбылоrS  X   принЯтьrT  X   прИнялrU  X   прИнялиrV  X   принялАrW  X   принУдитьrX  X
   рвАтьrY  X
   рвалАrZ  X   сверлИтьr[  X   сверлИшьr\  X   сверлИтr]  X
   снЯтьr^  X
   снялАr_  X   создАтьr`  X   создалАra  X   сорвАтьrb  X   сорвалАrc  X   сорИтьrd  X
   сорИтre  X   убрАтьrf  X   убралАrg  X   убыстрИтьrh  X   углубИтьri  X   укрепИтьrj  X   укрепИтrk  X   чЕрпатьrl  X   щемИтьrm  X
   щемИтrn  X   щЁлкатьro  X   балОванныйrp  X   включЁнныйrq  X   включЁнrr  X   низведЁнныйrs  X   довезЁнныйrt  X   зАгнутыйru  X   зАнятыйrv  X   занятАrw  X   зАпертыйrx  X   запертАry  X   заселЁнныйrz  X   заселенАr{  X   избалОванныйr|  X   балОванныйr}  X   кормЯщийr~  X   кровоточАщийr  X   молЯщийr�  X   нажИвшийr�  X   нАжитыйr�  X   нажитАr�  X   налИвшийr�  X   налитАr�  X   нанЯвшийся	r�  X   начАвшийr�  X   нАчатыйr�  X   низведЁнныйr�  X   низведЁнr�  X   включЁнныйr�  X   ободрЁнныйr�  X   ободрЁнr�  X   ободренАr�  X   обострЁнныйr�  X   отключЁнныйr�  X   определЁнныйr�  X   определЁнr�  X   отключЁнныйr�  X   повторЁнныйr�  X   поделЁнныйr�  X   понЯвшийr�  X   прИнятыйr�  X   приручЁнныйr�  X   прожИвшийr�  X   снЯтыйr�  X
   снятАr�  X   сОгнутыйr�  X   балУясьr�  X   закУпоривr�  X
   начАвr�  X   начАвшисьr�  X
   отдАвr�  X   поднЯвr�  X
   понЯвr�  X   прибЫвr�  X   вОвремяr�  X   добелАr�  X   дОверхуr�  X   донЕльзяr�  X   дОнизуr�  X   дОсухаr�  X   завИдноr�  X   зАгодяr�  X   зАсветлоr�  X   зАтемноr�  X   красИвееr�  X   навЕрхr�  X   надОлгоr�  X   ненадОлгоr�  e]r�  ej?  }r�  (jZ  ]r�  (KK K eX   лИтьсяr�  ]r�  (KK K ej�  ]r�  (K KKeuj\  j�  j]  ]r�  j�  aj_  ]r�  j�  aubJ牥;h)�r�  }r�  (h	J牥;h
X   Bahadirr�  hNh]r�  (]r�  ]r�  (j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  (j
  ]r�  (KK K ej  ]r�  (KK Kej  ]r�  (KK Keuj\  j�  j]  ]r�  j  aj_  ]r�  j  aubJ�(/h)�r�  }r�  (h	J�(/h
X   Dariar�  hNh]r�  (]r�  ]r�  (j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  (jY  ]r�  (KK K ej�  ]r�  (KK K ejf  ]r�  (KK K ej�  ]r�  (KK Kej�  ]r�  (KK K ej�  ]r�  (KK K ej�  ]r�  (KK K euj\  j*  j]  ]r�  j_  ]r�  ubJo(Bh)�r�  }r�  (h	Jo(Bh
X   🐊Простой🐊r�  hNh]r�  (]r�  ]r�  (j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j   j  j  j  j  j  j  j  j  j	  j
  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j   j!  j"  j#  j$  j%  j&  j'  j(  j)  j*  j+  j,  j-  j.  j/  j0  j1  j2  j3  j4  j5  j6  j7  j8  j9  j:  j;  j<  j=  j>  j?  j@  jA  jB  jC  jD  jE  jF  jG  jH  jI  jJ  jK  jL  jM  jN  jO  jP  jQ  jR  jS  jT  jU  jV  jW  jX  jY  jZ  j[  j\  j]  j^  j_  j`  ja  jb  jc  jd  je  jf  jg  jh  ji  jj  jk  jl  jm  jn  jo  jp  jq  jr  js  jt  ju  jv  jw  jx  jy  jz  j{  j|  j}  j~  j  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e]r�  ej?  }r�  j\  j�  j]  ]r�  j_  ]r�  ubu}r�  cbuiltins
set
r�  ]r�  �r�  Rr�  eX   periodr�  KX	   save_namer�  X   save.svr�  X   to_stopr�  �X   last_save_datetimer�  cdatetime
datetime
r�  C
�
(-�r�  �r�  Rr�  ub.